module aes (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire n_11512_o_0;
 wire n_11511_o_0;
 wire n_11510_o_0;
 wire n_11509_o_0;
 wire n_11508_o_0;
 wire _00410_;
 wire _00411_;
 wire n_11507_o_0;
 wire _00413_;
 wire n_11506_o_0;
 wire n_11505_o_0;
 wire n_11504_o_0;
 wire _00417_;
 wire n_11503_o_0;
 wire n_11502_o_0;
 wire n_11501_o_0;
 wire n_11500_o_0;
 wire n_11499_o_0;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire n_11498_o_0;
 wire n_11497_o_0;
 wire n_11496_o_0;
 wire n_11495_o_0;
 wire n_11494_o_0;
 wire n_11493_o_0;
 wire n_11492_o_0;
 wire n_11491_o_0;
 wire n_11490_o_0;
 wire n_11489_o_0;
 wire n_11488_o_0;
 wire n_11487_o_0;
 wire n_11486_o_0;
 wire n_11485_o_0;
 wire n_11484_o_0;
 wire n_11483_o_0;
 wire n_11482_o_0;
 wire n_11481_o_0;
 wire n_11480_o_0;
 wire n_11479_o_0;
 wire n_11478_o_0;
 wire n_11477_o_0;
 wire n_11476_o_0;
 wire n_11475_o_0;
 wire n_11474_o_0;
 wire n_11473_o_0;
 wire n_11472_o_0;
 wire n_11471_o_0;
 wire n_11470_o_0;
 wire n_11469_o_0;
 wire n_11468_o_0;
 wire n_11467_o_0;
 wire n_11466_o_0;
 wire n_11465_o_0;
 wire n_11464_o_0;
 wire _00489_;
 wire _00490_;
 wire n_11463_o_0;
 wire _00492_;
 wire n_11462_o_0;
 wire n_11461_o_0;
 wire n_11460_o_0;
 wire n_11459_o_0;
 wire n_11458_o_0;
 wire n_11457_o_0;
 wire _00499_;
 wire _00500_;
 wire n_11456_o_0;
 wire _00502_;
 wire n_11455_o_0;
 wire n_11454_o_0;
 wire n_11453_o_0;
 wire n_11452_o_0;
 wire n_11451_o_0;
 wire n_11450_o_0;
 wire _00509_;
 wire _00510_;
 wire n_11449_o_0;
 wire _00512_;
 wire n_11448_o_0;
 wire n_11447_o_0;
 wire n_11446_o_0;
 wire n_11445_o_0;
 wire n_11444_o_0;
 wire n_11443_o_0;
 wire _00519_;
 wire _00520_;
 wire n_11442_o_0;
 wire _00522_;
 wire n_11441_o_0;
 wire n_11440_o_0;
 wire n_11439_o_0;
 wire n_11438_o_0;
 wire n_11437_o_0;
 wire n_11436_o_0;
 wire _00529_;
 wire _00530_;
 wire n_11435_o_0;
 wire _00532_;
 wire n_11434_o_0;
 wire n_11433_o_0;
 wire n_11432_o_0;
 wire n_11431_o_0;
 wire n_11430_o_0;
 wire n_11429_o_0;
 wire _00539_;
 wire _00540_;
 wire n_11428_o_0;
 wire _00542_;
 wire n_11427_o_0;
 wire n_11426_o_0;
 wire n_11425_o_0;
 wire n_11424_o_0;
 wire n_11423_o_0;
 wire n_11422_o_0;
 wire _00549_;
 wire _00550_;
 wire n_11421_o_0;
 wire _00552_;
 wire n_11420_o_0;
 wire n_11419_o_0;
 wire n_11418_o_0;
 wire n_11417_o_0;
 wire n_11416_o_0;
 wire n_11415_o_0;
 wire _00559_;
 wire _00560_;
 wire n_11414_o_0;
 wire _00562_;
 wire n_11413_o_0;
 wire n_11412_o_0;
 wire n_11411_o_0;
 wire n_11410_o_0;
 wire n_11409_o_0;
 wire n_11408_o_0;
 wire _00569_;
 wire _00570_;
 wire n_11407_o_0;
 wire _00572_;
 wire n_11406_o_0;
 wire n_11405_o_0;
 wire n_11404_o_0;
 wire n_11403_o_0;
 wire n_11402_o_0;
 wire n_11401_o_0;
 wire n_11400_o_0;
 wire n_11399_o_0;
 wire _00581_;
 wire _00582_;
 wire n_11398_o_0;
 wire _00584_;
 wire n_11397_o_0;
 wire n_11396_o_0;
 wire n_11395_o_0;
 wire n_11394_o_0;
 wire n_11393_o_0;
 wire n_11392_o_0;
 wire n_11391_o_0;
 wire n_11390_o_0;
 wire _00593_;
 wire _00594_;
 wire n_11389_o_0;
 wire _00596_;
 wire n_11388_o_0;
 wire n_11387_o_0;
 wire n_11386_o_0;
 wire n_11385_o_0;
 wire n_11384_o_0;
 wire n_11383_o_0;
 wire n_11382_o_0;
 wire n_11381_o_0;
 wire _00605_;
 wire _00606_;
 wire n_11380_o_0;
 wire _00608_;
 wire n_11379_o_0;
 wire n_11378_o_0;
 wire n_11377_o_0;
 wire n_11376_o_0;
 wire n_11375_o_0;
 wire n_11374_o_0;
 wire n_11373_o_0;
 wire n_11372_o_0;
 wire _00617_;
 wire _00618_;
 wire n_11371_o_0;
 wire _00620_;
 wire n_11370_o_0;
 wire n_11369_o_0;
 wire n_11368_o_0;
 wire n_11367_o_0;
 wire n_11366_o_0;
 wire n_11365_o_0;
 wire _00627_;
 wire _00628_;
 wire n_11364_o_0;
 wire _00630_;
 wire n_11363_o_0;
 wire n_11362_o_0;
 wire n_11361_o_0;
 wire n_11360_o_0;
 wire n_11359_o_0;
 wire n_11358_o_0;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire n_11357_o_0;
 wire n_11356_o_0;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire n_11355_o_0;
 wire n_11354_o_0;
 wire n_11353_o_0;
 wire n_11352_o_0;
 wire n_11351_o_0;
 wire n_11350_o_0;
 wire n_11349_o_0;
 wire n_11348_o_0;
 wire n_11347_o_0;
 wire n_11346_o_0;
 wire n_11345_o_0;
 wire n_11344_o_0;
 wire n_11343_o_0;
 wire n_11342_o_0;
 wire n_11341_o_0;
 wire n_11340_o_0;
 wire n_11339_o_0;
 wire n_11338_o_0;
 wire n_11337_o_0;
 wire n_11336_o_0;
 wire n_11335_o_0;
 wire n_11334_o_0;
 wire n_11333_o_0;
 wire n_11332_o_0;
 wire n_11331_o_0;
 wire n_11330_o_0;
 wire n_11329_o_0;
 wire n_11328_o_0;
 wire n_11327_o_0;
 wire n_11326_o_0;
 wire n_11325_o_0;
 wire n_11324_o_0;
 wire n_11323_o_0;
 wire n_11322_o_0;
 wire n_11321_o_0;
 wire n_11320_o_0;
 wire n_11319_o_0;
 wire n_11318_o_0;
 wire n_11317_o_0;
 wire n_11316_o_0;
 wire n_11315_o_0;
 wire n_11314_o_0;
 wire n_11313_o_0;
 wire n_11312_o_0;
 wire n_11311_o_0;
 wire n_11310_o_0;
 wire n_11309_o_0;
 wire n_11308_o_0;
 wire n_11307_o_0;
 wire n_11306_o_0;
 wire n_11305_o_0;
 wire n_11304_o_0;
 wire n_11303_o_0;
 wire n_11302_o_0;
 wire n_11301_o_0;
 wire n_11300_o_0;
 wire n_11299_o_0;
 wire n_11298_o_0;
 wire n_11297_o_0;
 wire n_11296_o_0;
 wire n_11295_o_0;
 wire n_11294_o_0;
 wire n_11293_o_0;
 wire n_11292_o_0;
 wire n_11291_o_0;
 wire n_11290_o_0;
 wire n_11289_o_0;
 wire n_11288_o_0;
 wire n_11287_o_0;
 wire n_11286_o_0;
 wire n_11285_o_0;
 wire n_11284_o_0;
 wire n_11283_o_0;
 wire n_11282_o_0;
 wire n_11281_o_0;
 wire n_11280_o_0;
 wire n_11279_o_0;
 wire n_11278_o_0;
 wire n_11277_o_0;
 wire n_11276_o_0;
 wire n_11275_o_0;
 wire n_11274_o_0;
 wire n_11273_o_0;
 wire n_11272_o_0;
 wire n_11271_o_0;
 wire n_11270_o_0;
 wire n_11269_o_0;
 wire n_11268_o_0;
 wire n_11267_o_0;
 wire n_11266_o_0;
 wire n_11265_o_0;
 wire n_11264_o_0;
 wire n_11263_o_0;
 wire n_11262_o_0;
 wire n_11261_o_0;
 wire n_11260_o_0;
 wire n_11259_o_0;
 wire n_11258_o_0;
 wire n_11257_o_0;
 wire n_11256_o_0;
 wire n_11255_o_0;
 wire n_11254_o_0;
 wire n_11253_o_0;
 wire n_11252_o_0;
 wire n_11251_o_0;
 wire n_11250_o_0;
 wire n_11249_o_0;
 wire n_11248_o_0;
 wire n_11247_o_0;
 wire n_11246_o_0;
 wire n_11245_o_0;
 wire n_11244_o_0;
 wire n_11243_o_0;
 wire n_11242_o_0;
 wire n_11241_o_0;
 wire n_11240_o_0;
 wire n_11239_o_0;
 wire n_11238_o_0;
 wire n_11237_o_0;
 wire n_11236_o_0;
 wire n_11235_o_0;
 wire n_11234_o_0;
 wire n_11233_o_0;
 wire n_11232_o_0;
 wire n_11231_o_0;
 wire n_11230_o_0;
 wire n_11229_o_0;
 wire n_11228_o_0;
 wire n_11227_o_0;
 wire n_11226_o_0;
 wire n_11225_o_0;
 wire n_11224_o_0;
 wire n_11223_o_0;
 wire n_11222_o_0;
 wire n_11221_o_0;
 wire n_11220_o_0;
 wire n_11219_o_0;
 wire n_11218_o_0;
 wire n_11217_o_0;
 wire n_11216_o_0;
 wire n_11215_o_0;
 wire n_11214_o_0;
 wire n_11213_o_0;
 wire n_11212_o_0;
 wire n_11211_o_0;
 wire n_11210_o_0;
 wire n_11209_o_0;
 wire n_11208_o_0;
 wire n_11207_o_0;
 wire n_11206_o_0;
 wire n_11205_o_0;
 wire n_11204_o_0;
 wire n_11203_o_0;
 wire n_11202_o_0;
 wire n_11201_o_0;
 wire n_11200_o_0;
 wire n_11199_o_0;
 wire n_11198_o_0;
 wire n_11197_o_0;
 wire n_11196_o_0;
 wire n_11195_o_0;
 wire n_11194_o_0;
 wire n_11193_o_0;
 wire n_11192_o_0;
 wire n_11191_o_0;
 wire n_11190_o_0;
 wire n_11189_o_0;
 wire n_11188_o_0;
 wire n_11187_o_0;
 wire n_11186_o_0;
 wire n_11185_o_0;
 wire n_11184_o_0;
 wire n_11183_o_0;
 wire n_11182_o_0;
 wire n_11181_o_0;
 wire n_11180_o_0;
 wire n_11179_o_0;
 wire n_11178_o_0;
 wire n_11177_o_1;
 wire n_11177_o_0;
 wire n_11176_o_0;
 wire n_11175_o_0;
 wire n_11174_o_0;
 wire n_11173_o_0;
 wire n_11172_o_0;
 wire n_11171_o_0;
 wire n_11170_o_0;
 wire n_11169_o_0;
 wire n_11168_o_0;
 wire n_11167_o_0;
 wire n_11166_o_0;
 wire n_11165_o_0;
 wire n_11164_o_0;
 wire n_11163_o_0;
 wire n_11162_o_0;
 wire n_11161_o_0;
 wire n_11160_o_0;
 wire n_11159_o_0;
 wire n_11158_o_0;
 wire n_11157_o_0;
 wire n_11156_o_0;
 wire n_11155_o_0;
 wire n_11154_o_0;
 wire n_11153_o_0;
 wire n_11152_o_0;
 wire n_11151_o_0;
 wire n_11150_o_0;
 wire n_11149_o_0;
 wire n_11148_o_0;
 wire n_11147_o_0;
 wire n_11146_o_0;
 wire n_11145_o_0;
 wire n_11144_o_0;
 wire n_11143_o_0;
 wire n_11142_o_0;
 wire n_11141_o_0;
 wire n_11140_o_0;
 wire n_11139_o_0;
 wire n_11138_o_0;
 wire n_11137_o_0;
 wire n_11136_o_0;
 wire n_11135_o_0;
 wire n_11134_o_0;
 wire n_11133_o_0;
 wire n_11132_o_0;
 wire n_11131_o_0;
 wire n_11130_o_0;
 wire n_11129_o_0;
 wire n_11128_o_0;
 wire n_11127_o_0;
 wire n_11126_o_0;
 wire n_11125_o_0;
 wire n_11124_o_0;
 wire n_11123_o_0;
 wire n_11122_o_0;
 wire n_11121_o_0;
 wire n_11120_o_0;
 wire n_11119_o_0;
 wire n_11118_o_0;
 wire n_11117_o_0;
 wire n_11116_o_0;
 wire n_11115_o_0;
 wire n_11114_o_0;
 wire n_11113_o_0;
 wire n_11112_o_0;
 wire n_11111_o_0;
 wire n_11110_o_0;
 wire n_11109_o_0;
 wire n_11108_o_0;
 wire n_11107_o_0;
 wire n_11106_o_0;
 wire n_11105_o_0;
 wire n_11104_o_0;
 wire n_11103_o_0;
 wire n_11102_o_0;
 wire n_11101_o_0;
 wire n_11100_o_0;
 wire n_11099_o_0;
 wire n_11098_o_0;
 wire n_11097_o_0;
 wire n_11096_o_0;
 wire n_11095_o_0;
 wire n_11094_o_0;
 wire n_11093_o_0;
 wire n_11092_o_0;
 wire n_11091_o_0;
 wire n_11090_o_0;
 wire n_11089_o_0;
 wire n_11088_o_0;
 wire n_11087_o_0;
 wire n_11086_o_0;
 wire n_11085_o_0;
 wire n_11084_o_0;
 wire n_11083_o_0;
 wire n_11082_o_0;
 wire n_11081_o_0;
 wire n_11080_o_0;
 wire n_11079_o_0;
 wire n_11078_o_0;
 wire n_11077_o_0;
 wire n_11076_o_0;
 wire n_11075_o_0;
 wire n_11074_o_0;
 wire n_11073_o_0;
 wire n_11072_o_0;
 wire n_11071_o_0;
 wire n_11070_o_0;
 wire n_11069_o_0;
 wire n_11068_o_0;
 wire n_11067_o_0;
 wire n_11066_o_0;
 wire n_11065_o_0;
 wire n_11064_o_0;
 wire n_11063_o_0;
 wire n_11062_o_0;
 wire n_11061_o_0;
 wire n_11060_o_0;
 wire n_11059_o_0;
 wire n_11058_o_0;
 wire n_11057_o_0;
 wire n_11056_o_0;
 wire n_11055_o_0;
 wire n_11054_o_0;
 wire n_11053_o_0;
 wire n_11052_o_0;
 wire n_11051_o_0;
 wire n_11050_o_0;
 wire n_11049_o_0;
 wire n_11048_o_0;
 wire n_11047_o_0;
 wire n_11046_o_0;
 wire n_11045_o_0;
 wire n_11044_o_0;
 wire n_11043_o_0;
 wire n_11042_o_0;
 wire n_11041_o_0;
 wire n_11040_o_0;
 wire n_11039_o_0;
 wire n_11038_o_0;
 wire n_11037_o_0;
 wire n_11036_o_0;
 wire n_11035_o_0;
 wire n_11034_o_0;
 wire n_11033_o_0;
 wire n_11032_o_0;
 wire n_11031_o_0;
 wire n_11030_o_0;
 wire n_11029_o_0;
 wire n_11028_o_0;
 wire n_11027_o_0;
 wire n_11026_o_0;
 wire n_11025_o_0;
 wire n_11024_o_0;
 wire n_11023_o_0;
 wire n_11022_o_0;
 wire n_11021_o_0;
 wire n_11020_o_0;
 wire n_11019_o_0;
 wire n_11018_o_0;
 wire n_11017_o_0;
 wire n_11016_o_0;
 wire n_11015_o_0;
 wire n_11014_o_0;
 wire n_11013_o_0;
 wire n_11012_o_0;
 wire n_11011_o_0;
 wire n_11010_o_0;
 wire n_11009_o_0;
 wire n_11008_o_0;
 wire n_11007_o_0;
 wire n_11006_o_0;
 wire n_11005_o_0;
 wire n_11004_o_0;
 wire n_11003_o_0;
 wire n_11002_o_0;
 wire n_11001_o_0;
 wire n_11000_o_0;
 wire n_10999_o_0;
 wire n_10998_o_0;
 wire n_10997_o_0;
 wire n_10996_o_0;
 wire n_10995_o_0;
 wire n_10994_o_0;
 wire n_10993_o_0;
 wire n_10992_o_0;
 wire n_10991_o_0;
 wire n_10990_o_0;
 wire n_10989_o_0;
 wire n_10988_o_0;
 wire n_10987_o_0;
 wire n_10986_o_0;
 wire n_10985_o_0;
 wire n_10984_o_0;
 wire n_10983_o_0;
 wire n_10982_o_0;
 wire n_10981_o_0;
 wire n_10980_o_0;
 wire n_10979_o_0;
 wire n_10978_o_0;
 wire n_10977_o_0;
 wire n_10976_o_0;
 wire n_10975_o_0;
 wire n_10974_o_0;
 wire n_10973_o_0;
 wire n_10972_o_0;
 wire n_10971_o_0;
 wire n_10970_o_0;
 wire n_10969_o_0;
 wire n_10968_o_0;
 wire n_10967_o_0;
 wire n_10966_o_0;
 wire n_10965_o_0;
 wire n_10964_o_0;
 wire n_10963_o_0;
 wire n_10962_o_0;
 wire n_10961_o_0;
 wire n_10960_o_0;
 wire n_10959_o_0;
 wire n_10958_o_0;
 wire n_10957_o_0;
 wire n_10956_o_0;
 wire n_10955_o_0;
 wire n_10954_o_0;
 wire n_10953_o_0;
 wire n_10952_o_0;
 wire n_10951_o_0;
 wire n_10950_o_0;
 wire n_10949_o_0;
 wire n_10948_o_0;
 wire n_10947_o_0;
 wire n_10946_o_0;
 wire n_10945_o_0;
 wire n_10944_o_0;
 wire n_10943_o_0;
 wire n_10942_o_0;
 wire n_10941_o_0;
 wire n_10940_o_0;
 wire n_10939_o_0;
 wire n_10938_o_0;
 wire n_10937_o_0;
 wire n_10936_o_0;
 wire n_10935_o_0;
 wire n_10934_o_0;
 wire n_10933_o_0;
 wire n_10932_o_0;
 wire n_10931_o_0;
 wire n_10930_o_0;
 wire n_10929_o_0;
 wire n_10928_o_0;
 wire n_10927_o_0;
 wire n_10926_o_0;
 wire n_10925_o_0;
 wire n_10924_o_0;
 wire n_10923_o_0;
 wire n_10922_o_0;
 wire n_10921_o_0;
 wire n_10920_o_0;
 wire n_10919_o_0;
 wire n_10918_o_0;
 wire n_10917_o_0;
 wire n_10916_o_0;
 wire n_10915_o_0;
 wire n_10914_o_0;
 wire n_10913_o_0;
 wire n_10912_o_0;
 wire n_10911_o_0;
 wire n_10910_o_0;
 wire n_10909_o_0;
 wire n_10908_o_0;
 wire n_10907_o_0;
 wire n_10906_o_0;
 wire n_10905_o_0;
 wire n_10904_o_0;
 wire n_10903_o_0;
 wire n_10902_o_0;
 wire n_10901_o_0;
 wire n_10900_o_0;
 wire n_10899_o_0;
 wire n_10898_o_0;
 wire n_10897_o_0;
 wire n_10896_o_0;
 wire n_10895_o_0;
 wire n_10894_o_0;
 wire n_10893_o_0;
 wire n_10892_o_0;
 wire n_10891_o_0;
 wire n_10890_o_0;
 wire n_10889_o_0;
 wire n_10888_o_0;
 wire n_10887_o_0;
 wire n_10886_o_0;
 wire n_10885_o_0;
 wire n_10884_o_0;
 wire n_10883_o_0;
 wire n_10882_o_0;
 wire n_10881_o_0;
 wire n_10880_o_0;
 wire n_10879_o_0;
 wire n_10878_o_0;
 wire n_10877_o_0;
 wire n_10876_o_0;
 wire n_10875_o_0;
 wire n_10874_o_0;
 wire n_10873_o_0;
 wire n_10872_o_0;
 wire n_10871_o_0;
 wire n_10870_o_0;
 wire n_10869_o_0;
 wire n_10868_o_0;
 wire n_10867_o_0;
 wire n_10866_o_0;
 wire n_10865_o_0;
 wire n_10864_o_0;
 wire n_10863_o_0;
 wire n_10862_o_0;
 wire n_10861_o_0;
 wire n_10860_o_0;
 wire n_10859_o_0;
 wire n_10858_o_0;
 wire n_10857_o_0;
 wire n_10856_o_0;
 wire n_10855_o_0;
 wire n_10854_o_0;
 wire n_10853_o_0;
 wire n_10852_o_0;
 wire n_10851_o_0;
 wire n_10850_o_0;
 wire n_10849_o_0;
 wire n_10848_o_0;
 wire n_10847_o_0;
 wire n_10846_o_0;
 wire n_10845_o_0;
 wire n_10844_o_0;
 wire n_10843_o_0;
 wire n_10842_o_0;
 wire n_10841_o_0;
 wire n_10840_o_0;
 wire n_10839_o_0;
 wire n_10838_o_0;
 wire n_10837_o_0;
 wire n_10836_o_0;
 wire n_10835_o_0;
 wire n_10834_o_0;
 wire n_10833_o_0;
 wire n_10832_o_0;
 wire n_10831_o_0;
 wire n_10830_o_0;
 wire n_10829_o_0;
 wire n_10828_o_0;
 wire n_10827_o_0;
 wire n_10826_o_0;
 wire n_10825_o_0;
 wire n_10824_o_0;
 wire n_10823_o_0;
 wire n_10822_o_0;
 wire n_10821_o_0;
 wire n_10820_o_0;
 wire n_10819_o_0;
 wire n_10818_o_0;
 wire n_10817_o_0;
 wire n_10816_o_0;
 wire n_10815_o_0;
 wire n_10814_o_0;
 wire n_10813_o_0;
 wire n_10812_o_0;
 wire n_10811_o_0;
 wire n_10810_o_0;
 wire n_10809_o_0;
 wire n_10808_o_0;
 wire n_10807_o_0;
 wire n_10806_o_0;
 wire n_10805_o_0;
 wire n_10804_o_0;
 wire n_10803_o_0;
 wire n_10802_o_0;
 wire n_10801_o_0;
 wire n_10800_o_0;
 wire n_10799_o_0;
 wire n_10798_o_0;
 wire n_10797_o_0;
 wire n_10796_o_0;
 wire n_10795_o_0;
 wire n_10794_o_0;
 wire n_10793_o_0;
 wire n_10792_o_0;
 wire n_10791_o_0;
 wire n_10790_o_0;
 wire n_10789_o_0;
 wire n_10788_o_0;
 wire n_10787_o_0;
 wire n_10786_o_0;
 wire n_10785_o_0;
 wire n_10784_o_0;
 wire n_10783_o_0;
 wire n_10782_o_0;
 wire n_10781_o_0;
 wire n_10780_o_0;
 wire n_10779_o_0;
 wire n_10778_o_0;
 wire n_10777_o_0;
 wire n_10776_o_0;
 wire n_10775_o_0;
 wire n_10774_o_0;
 wire n_10773_o_0;
 wire n_10772_o_0;
 wire n_10771_o_0;
 wire n_10770_o_0;
 wire n_10769_o_0;
 wire n_10768_o_0;
 wire n_10767_o_0;
 wire n_10766_o_0;
 wire n_10765_o_0;
 wire n_10764_o_0;
 wire n_10763_o_0;
 wire n_10762_o_0;
 wire n_10761_o_0;
 wire n_10760_o_0;
 wire n_10759_o_0;
 wire n_10758_o_0;
 wire n_10757_o_0;
 wire n_10756_o_0;
 wire n_10755_o_0;
 wire n_10754_o_0;
 wire n_10753_o_0;
 wire n_10752_o_0;
 wire n_10751_o_0;
 wire n_10750_o_0;
 wire n_10749_o_0;
 wire n_10748_o_0;
 wire n_10747_o_0;
 wire n_10746_o_0;
 wire n_10745_o_0;
 wire n_10744_o_0;
 wire n_10743_o_0;
 wire n_10742_o_0;
 wire n_10741_o_0;
 wire n_10740_o_0;
 wire n_10739_o_0;
 wire n_10738_o_0;
 wire n_10737_o_0;
 wire n_10736_o_0;
 wire n_10735_o_0;
 wire n_10734_o_0;
 wire n_10733_o_0;
 wire n_10732_o_0;
 wire n_10731_o_0;
 wire n_10730_o_0;
 wire n_10729_o_0;
 wire n_10728_o_0;
 wire n_10727_o_0;
 wire n_10726_o_0;
 wire n_10725_o_0;
 wire n_10724_o_0;
 wire n_10723_o_0;
 wire n_10722_o_0;
 wire n_10721_o_0;
 wire n_10720_o_0;
 wire n_10719_o_0;
 wire n_10718_o_0;
 wire n_10717_o_0;
 wire n_10716_o_0;
 wire n_10715_o_0;
 wire n_10714_o_0;
 wire n_10713_o_0;
 wire n_10712_o_0;
 wire n_10711_o_0;
 wire n_10710_o_0;
 wire n_10709_o_0;
 wire n_10708_o_0;
 wire n_10707_o_0;
 wire n_10706_o_0;
 wire n_10705_o_0;
 wire n_10704_o_0;
 wire n_10703_o_0;
 wire n_10702_o_0;
 wire n_10701_o_0;
 wire n_10700_o_0;
 wire n_10699_o_0;
 wire n_10698_o_0;
 wire n_10697_o_0;
 wire n_10696_o_0;
 wire n_10695_o_0;
 wire n_10694_o_0;
 wire n_10693_o_0;
 wire n_10692_o_0;
 wire n_10691_o_0;
 wire n_10690_o_0;
 wire n_10689_o_0;
 wire n_10688_o_0;
 wire n_10687_o_0;
 wire n_10686_o_0;
 wire n_10685_o_0;
 wire n_10684_o_0;
 wire n_10683_o_0;
 wire n_10682_o_0;
 wire n_10681_o_0;
 wire n_10680_o_0;
 wire n_10679_o_0;
 wire n_10678_o_0;
 wire n_10677_o_0;
 wire n_10676_o_0;
 wire n_10675_o_0;
 wire n_10674_o_0;
 wire n_10673_o_0;
 wire n_10672_o_0;
 wire n_10671_o_0;
 wire n_10670_o_0;
 wire n_10669_o_0;
 wire n_10668_o_0;
 wire n_10667_o_0;
 wire n_10666_o_0;
 wire n_10665_o_0;
 wire n_10664_o_0;
 wire n_10663_o_0;
 wire n_10662_o_0;
 wire n_10661_o_0;
 wire n_10660_o_0;
 wire n_10659_o_0;
 wire n_10658_o_0;
 wire n_10657_o_0;
 wire n_10656_o_0;
 wire n_10655_o_0;
 wire n_10654_o_0;
 wire n_10653_o_0;
 wire n_10652_o_0;
 wire n_10651_o_0;
 wire n_10650_o_0;
 wire n_10649_o_0;
 wire n_10648_o_0;
 wire n_10647_o_0;
 wire n_10646_o_0;
 wire n_10645_o_0;
 wire n_10644_o_0;
 wire n_10643_o_0;
 wire n_10642_o_0;
 wire n_10641_o_0;
 wire n_10640_o_0;
 wire n_10639_o_0;
 wire n_10638_o_0;
 wire n_10637_o_0;
 wire n_10636_o_0;
 wire n_10635_o_0;
 wire n_10634_o_0;
 wire n_10633_o_0;
 wire n_10632_o_0;
 wire n_10631_o_0;
 wire n_10630_o_0;
 wire n_10629_o_0;
 wire n_10628_o_0;
 wire n_10627_o_0;
 wire n_10626_o_0;
 wire n_10625_o_0;
 wire n_10624_o_0;
 wire n_10623_o_0;
 wire n_10622_o_0;
 wire n_10621_o_0;
 wire n_10620_o_0;
 wire n_10619_o_0;
 wire n_10618_o_0;
 wire n_10617_o_0;
 wire n_10616_o_0;
 wire n_10615_o_0;
 wire n_10614_o_0;
 wire n_10613_o_0;
 wire n_10612_o_0;
 wire n_10611_o_0;
 wire n_10610_o_0;
 wire n_10609_o_0;
 wire n_10608_o_0;
 wire n_10607_o_0;
 wire n_10606_o_0;
 wire n_10605_o_0;
 wire n_10604_o_0;
 wire n_10603_o_0;
 wire n_10602_o_0;
 wire n_10601_o_0;
 wire n_10600_o_0;
 wire n_10599_o_0;
 wire n_10598_o_0;
 wire n_10597_o_0;
 wire n_10596_o_0;
 wire n_10595_o_0;
 wire n_10594_o_0;
 wire n_10593_o_0;
 wire n_10592_o_0;
 wire n_10591_o_0;
 wire n_10590_o_0;
 wire n_10589_o_0;
 wire n_10588_o_0;
 wire n_10587_o_0;
 wire n_10586_o_0;
 wire n_10585_o_0;
 wire n_10584_o_0;
 wire n_10583_o_0;
 wire n_10582_o_0;
 wire n_10581_o_0;
 wire n_10580_o_0;
 wire n_10579_o_0;
 wire n_10578_o_0;
 wire n_10577_o_0;
 wire n_10576_o_0;
 wire n_10575_o_0;
 wire n_10574_o_0;
 wire n_10573_o_0;
 wire n_10572_o_0;
 wire n_10571_o_0;
 wire n_10570_o_0;
 wire n_10569_o_0;
 wire n_10568_o_0;
 wire n_10567_o_0;
 wire n_10566_o_0;
 wire n_10565_o_0;
 wire n_10564_o_0;
 wire n_10563_o_0;
 wire n_10562_o_0;
 wire n_10561_o_0;
 wire n_10560_o_0;
 wire n_10559_o_0;
 wire n_10558_o_0;
 wire n_10557_o_0;
 wire n_10556_o_0;
 wire n_10555_o_0;
 wire n_10554_o_0;
 wire n_10553_o_0;
 wire n_10552_o_0;
 wire n_10551_o_0;
 wire n_10550_o_0;
 wire n_10549_o_0;
 wire n_10548_o_0;
 wire n_10547_o_0;
 wire n_10546_o_0;
 wire n_10545_o_0;
 wire n_10544_o_0;
 wire n_10543_o_0;
 wire n_10542_o_0;
 wire n_10541_o_0;
 wire n_10540_o_0;
 wire n_10539_o_0;
 wire n_10538_o_0;
 wire n_10537_o_0;
 wire n_10536_o_0;
 wire n_10535_o_0;
 wire n_10534_o_0;
 wire n_10533_o_0;
 wire n_10532_o_0;
 wire n_10531_o_0;
 wire n_10530_o_0;
 wire n_10529_o_0;
 wire n_10528_o_0;
 wire n_10527_o_0;
 wire n_10526_o_0;
 wire n_10525_o_0;
 wire n_10524_o_0;
 wire n_10523_o_0;
 wire n_10522_o_0;
 wire n_10521_o_0;
 wire n_10520_o_0;
 wire n_10519_o_0;
 wire n_10518_o_0;
 wire n_10517_o_0;
 wire n_10516_o_0;
 wire n_10515_o_0;
 wire n_10514_o_0;
 wire n_10513_o_0;
 wire n_10512_o_0;
 wire n_10511_o_0;
 wire n_10510_o_0;
 wire n_10509_o_0;
 wire n_10508_o_0;
 wire n_10507_o_0;
 wire n_10506_o_0;
 wire n_10505_o_0;
 wire n_10504_o_0;
 wire n_10503_o_0;
 wire n_10502_o_0;
 wire n_10501_o_0;
 wire n_10500_o_0;
 wire n_10499_o_0;
 wire n_10498_o_0;
 wire n_10497_o_0;
 wire n_10496_o_0;
 wire n_10495_o_0;
 wire n_10494_o_0;
 wire n_10493_o_0;
 wire n_10492_o_0;
 wire n_10491_o_0;
 wire n_10490_o_0;
 wire n_10489_o_0;
 wire n_10488_o_0;
 wire n_10487_o_0;
 wire n_10486_o_0;
 wire n_10485_o_0;
 wire n_10484_o_0;
 wire n_10483_o_0;
 wire n_10482_o_0;
 wire n_10481_o_0;
 wire n_10480_o_0;
 wire n_10479_o_0;
 wire n_10478_o_0;
 wire n_10477_o_0;
 wire n_10476_o_0;
 wire n_10475_o_0;
 wire n_10474_o_0;
 wire n_10473_o_0;
 wire n_10472_o_0;
 wire n_10471_o_0;
 wire n_10470_o_0;
 wire n_10469_o_0;
 wire n_10468_o_0;
 wire n_10467_o_0;
 wire n_10466_o_0;
 wire n_10465_o_0;
 wire n_10464_o_0;
 wire n_10463_o_0;
 wire n_10462_o_0;
 wire n_10461_o_0;
 wire n_10460_o_0;
 wire n_10459_o_0;
 wire n_10458_o_0;
 wire n_10457_o_0;
 wire n_10456_o_0;
 wire n_10455_o_0;
 wire n_10454_o_0;
 wire n_10453_o_0;
 wire n_10452_o_0;
 wire n_10451_o_0;
 wire n_10450_o_0;
 wire n_10449_o_0;
 wire n_10448_o_0;
 wire n_10447_o_0;
 wire n_10446_o_0;
 wire n_10445_o_0;
 wire n_10444_o_0;
 wire n_10443_o_0;
 wire n_10442_o_0;
 wire n_10441_o_0;
 wire n_10440_o_0;
 wire n_10439_o_0;
 wire n_10438_o_0;
 wire n_10437_o_0;
 wire n_10436_o_0;
 wire n_10435_o_0;
 wire n_10434_o_0;
 wire n_10433_o_0;
 wire n_10432_o_0;
 wire n_10431_o_0;
 wire n_10430_o_0;
 wire n_10429_o_0;
 wire n_10428_o_0;
 wire n_10427_o_0;
 wire n_10426_o_0;
 wire n_10425_o_0;
 wire n_10424_o_0;
 wire n_10423_o_0;
 wire n_10422_o_0;
 wire n_10421_o_0;
 wire n_10420_o_0;
 wire n_10419_o_0;
 wire n_10418_o_0;
 wire n_10417_o_0;
 wire n_10416_o_0;
 wire n_10415_o_0;
 wire n_10414_o_0;
 wire n_10413_o_0;
 wire n_10412_o_0;
 wire n_10411_o_0;
 wire n_10410_o_0;
 wire n_10409_o_0;
 wire n_10408_o_0;
 wire n_10407_o_0;
 wire n_10406_o_0;
 wire n_10405_o_0;
 wire n_10404_o_0;
 wire n_10403_o_0;
 wire n_10402_o_0;
 wire n_10401_o_0;
 wire n_10400_o_0;
 wire n_10399_o_0;
 wire n_10398_o_0;
 wire n_10397_o_0;
 wire n_10396_o_0;
 wire n_10395_o_0;
 wire n_10394_o_0;
 wire n_10393_o_0;
 wire n_10392_o_0;
 wire n_10391_o_0;
 wire n_10390_o_0;
 wire n_10389_o_0;
 wire n_10388_o_0;
 wire n_10387_o_0;
 wire n_10386_o_0;
 wire n_10385_o_0;
 wire n_10384_o_0;
 wire n_10383_o_0;
 wire n_10382_o_0;
 wire n_10381_o_0;
 wire n_10380_o_0;
 wire n_10379_o_0;
 wire n_10378_o_0;
 wire n_10377_o_0;
 wire n_10376_o_0;
 wire n_10375_o_0;
 wire n_10374_o_0;
 wire n_10373_o_0;
 wire n_10372_o_0;
 wire n_10371_o_0;
 wire n_10370_o_0;
 wire n_10369_o_0;
 wire n_10368_o_0;
 wire n_10367_o_0;
 wire n_10366_o_0;
 wire n_10365_o_0;
 wire n_10364_o_0;
 wire n_10363_o_0;
 wire n_10362_o_0;
 wire n_10361_o_0;
 wire n_10360_o_0;
 wire n_10359_o_0;
 wire n_10358_o_0;
 wire n_10357_o_0;
 wire n_10356_o_0;
 wire n_10355_o_0;
 wire n_10354_o_0;
 wire n_10353_o_0;
 wire n_10352_o_0;
 wire n_10351_o_0;
 wire n_10350_o_0;
 wire n_10349_o_0;
 wire n_10348_o_0;
 wire n_10347_o_0;
 wire n_10346_o_0;
 wire n_10345_o_0;
 wire n_10344_o_0;
 wire n_10343_o_0;
 wire n_10342_o_0;
 wire n_10341_o_0;
 wire n_10340_o_0;
 wire n_10339_o_0;
 wire n_10338_o_0;
 wire n_10337_o_0;
 wire n_10336_o_0;
 wire n_10335_o_0;
 wire n_10334_o_0;
 wire n_10333_o_0;
 wire n_10332_o_0;
 wire n_10331_o_0;
 wire n_10330_o_0;
 wire n_10329_o_0;
 wire n_10328_o_0;
 wire n_10327_o_0;
 wire n_10326_o_0;
 wire n_10325_o_0;
 wire n_10324_o_0;
 wire n_10323_o_0;
 wire n_10322_o_0;
 wire n_10321_o_0;
 wire n_10320_o_0;
 wire n_10319_o_0;
 wire n_10318_o_0;
 wire n_10317_o_0;
 wire n_10316_o_0;
 wire n_10315_o_0;
 wire n_10314_o_0;
 wire n_10313_o_0;
 wire n_10312_o_0;
 wire n_10311_o_0;
 wire n_10310_o_0;
 wire n_10309_o_0;
 wire n_10308_o_0;
 wire n_10307_o_0;
 wire n_10306_o_0;
 wire n_10305_o_0;
 wire n_10304_o_0;
 wire n_10303_o_0;
 wire n_10302_o_0;
 wire n_10301_o_0;
 wire n_10300_o_0;
 wire n_10299_o_0;
 wire n_10298_o_0;
 wire n_10297_o_0;
 wire n_10296_o_0;
 wire n_10295_o_0;
 wire n_10294_o_0;
 wire n_10293_o_0;
 wire n_10292_o_0;
 wire n_10291_o_0;
 wire n_10290_o_0;
 wire n_10289_o_0;
 wire n_10288_o_0;
 wire n_10287_o_0;
 wire n_10286_o_0;
 wire n_10285_o_0;
 wire n_10284_o_0;
 wire n_10283_o_0;
 wire n_10282_o_0;
 wire n_10281_o_0;
 wire n_10280_o_0;
 wire n_10279_o_0;
 wire n_10278_o_0;
 wire n_10277_o_0;
 wire n_10276_o_0;
 wire n_10275_o_0;
 wire n_10274_o_0;
 wire n_10273_o_0;
 wire n_10272_o_0;
 wire n_10271_o_0;
 wire n_10270_o_0;
 wire n_10269_o_0;
 wire n_10268_o_0;
 wire n_10267_o_0;
 wire n_10266_o_0;
 wire n_10265_o_0;
 wire n_10264_o_0;
 wire n_10263_o_0;
 wire n_10262_o_0;
 wire n_10261_o_0;
 wire n_10260_o_0;
 wire n_10259_o_0;
 wire n_10258_o_0;
 wire n_10257_o_0;
 wire n_10256_o_0;
 wire n_10255_o_0;
 wire n_10254_o_0;
 wire n_10253_o_0;
 wire n_10252_o_0;
 wire n_10251_o_0;
 wire n_10250_o_0;
 wire n_10249_o_0;
 wire n_10248_o_0;
 wire n_10247_o_0;
 wire n_10246_o_0;
 wire n_10245_o_0;
 wire n_10244_o_0;
 wire n_10243_o_0;
 wire n_10242_o_0;
 wire n_10241_o_0;
 wire n_10240_o_0;
 wire n_10239_o_0;
 wire n_10238_o_0;
 wire n_10237_o_0;
 wire n_10236_o_0;
 wire n_10235_o_0;
 wire n_10234_o_0;
 wire n_10233_o_0;
 wire n_10232_o_0;
 wire n_10231_o_0;
 wire n_10230_o_0;
 wire n_10229_o_0;
 wire n_10228_o_0;
 wire n_10227_o_0;
 wire n_10226_o_0;
 wire n_10225_o_0;
 wire n_10224_o_0;
 wire n_10223_o_0;
 wire n_10222_o_0;
 wire n_10221_o_0;
 wire n_10220_o_0;
 wire n_10219_o_0;
 wire n_10218_o_0;
 wire n_10217_o_0;
 wire n_10216_o_0;
 wire n_10215_o_0;
 wire n_10214_o_0;
 wire n_10213_o_0;
 wire n_10212_o_0;
 wire n_10211_o_0;
 wire n_10210_o_0;
 wire n_10209_o_0;
 wire n_10208_o_0;
 wire n_10207_o_0;
 wire n_10206_o_0;
 wire n_10205_o_0;
 wire n_10204_o_0;
 wire n_10203_o_0;
 wire n_10202_o_0;
 wire n_10201_o_0;
 wire n_10200_o_0;
 wire n_10199_o_0;
 wire n_10198_o_0;
 wire n_10197_o_0;
 wire n_10196_o_0;
 wire n_10195_o_0;
 wire n_10194_o_0;
 wire n_10193_o_0;
 wire n_10192_o_0;
 wire n_10191_o_0;
 wire n_10190_o_0;
 wire n_10189_o_0;
 wire n_10188_o_0;
 wire n_10187_o_0;
 wire n_10186_o_0;
 wire n_10185_o_0;
 wire n_10184_o_0;
 wire n_10183_o_0;
 wire n_10182_o_0;
 wire n_10181_o_0;
 wire n_10180_o_0;
 wire n_10179_o_0;
 wire n_10178_o_0;
 wire n_10177_o_0;
 wire n_10176_o_0;
 wire n_10175_o_0;
 wire n_10174_o_0;
 wire n_10173_o_0;
 wire n_10172_o_0;
 wire n_10171_o_0;
 wire n_10170_o_0;
 wire n_10169_o_0;
 wire n_10168_o_0;
 wire n_10167_o_0;
 wire n_10166_o_0;
 wire n_10165_o_0;
 wire n_10164_o_0;
 wire n_10163_o_0;
 wire n_10162_o_0;
 wire n_10161_o_0;
 wire n_10160_o_0;
 wire n_10159_o_0;
 wire n_10158_o_0;
 wire n_10157_o_0;
 wire n_10156_o_0;
 wire n_10155_o_0;
 wire n_10154_o_0;
 wire n_10153_o_0;
 wire n_10152_o_0;
 wire n_10151_o_0;
 wire n_10150_o_0;
 wire n_10149_o_0;
 wire n_10148_o_0;
 wire n_10147_o_0;
 wire n_10146_o_0;
 wire n_10145_o_0;
 wire n_10144_o_0;
 wire n_10143_o_0;
 wire n_10142_o_0;
 wire n_10141_o_0;
 wire n_10140_o_0;
 wire n_10139_o_0;
 wire n_10138_o_0;
 wire n_10137_o_0;
 wire n_10136_o_0;
 wire n_10135_o_0;
 wire n_10134_o_0;
 wire n_10133_o_0;
 wire n_10132_o_0;
 wire n_10131_o_0;
 wire n_10130_o_0;
 wire n_10129_o_0;
 wire n_10128_o_0;
 wire n_10127_o_0;
 wire n_10126_o_0;
 wire n_10125_o_0;
 wire n_10124_o_0;
 wire n_10123_o_0;
 wire n_10122_o_0;
 wire n_10121_o_0;
 wire n_10120_o_0;
 wire n_10119_o_0;
 wire n_10118_o_0;
 wire n_10117_o_0;
 wire n_10116_o_0;
 wire n_10115_o_0;
 wire n_10114_o_0;
 wire n_10113_o_0;
 wire n_10112_o_0;
 wire n_10111_o_0;
 wire n_10110_o_0;
 wire n_10109_o_0;
 wire n_10108_o_0;
 wire n_10107_o_0;
 wire n_10106_o_0;
 wire n_10105_o_0;
 wire n_10104_o_0;
 wire n_10103_o_0;
 wire n_10102_o_0;
 wire n_10101_o_0;
 wire n_10100_o_0;
 wire n_10099_o_0;
 wire n_10098_o_0;
 wire n_10097_o_0;
 wire n_10096_o_0;
 wire n_10095_o_0;
 wire n_10094_o_0;
 wire n_10093_o_0;
 wire n_10092_o_0;
 wire n_10091_o_0;
 wire n_10090_o_0;
 wire n_10089_o_0;
 wire n_10088_o_0;
 wire n_10087_o_0;
 wire n_10086_o_0;
 wire n_10085_o_0;
 wire n_10084_o_0;
 wire n_10083_o_0;
 wire n_10082_o_0;
 wire n_10081_o_0;
 wire n_10080_o_0;
 wire n_10079_o_0;
 wire n_10078_o_0;
 wire n_10077_o_0;
 wire n_10076_o_0;
 wire n_10075_o_0;
 wire n_10074_o_0;
 wire n_10073_o_0;
 wire n_10072_o_0;
 wire n_10071_o_0;
 wire n_10070_o_0;
 wire n_10069_o_0;
 wire n_10068_o_0;
 wire n_10067_o_0;
 wire n_10066_o_0;
 wire n_10065_o_0;
 wire n_10064_o_0;
 wire n_10063_o_0;
 wire n_10062_o_0;
 wire n_10061_o_0;
 wire n_10060_o_0;
 wire n_10059_o_0;
 wire n_10058_o_0;
 wire n_10057_o_0;
 wire n_10056_o_0;
 wire n_10055_o_0;
 wire n_10054_o_0;
 wire n_10053_o_0;
 wire n_10052_o_0;
 wire n_10051_o_0;
 wire n_10050_o_0;
 wire n_10049_o_0;
 wire n_10048_o_0;
 wire n_10047_o_0;
 wire n_10046_o_0;
 wire n_10045_o_0;
 wire n_10044_o_0;
 wire n_10043_o_0;
 wire n_10042_o_0;
 wire n_10041_o_0;
 wire n_10040_o_0;
 wire n_10039_o_0;
 wire n_10038_o_0;
 wire n_10037_o_0;
 wire n_10036_o_0;
 wire n_10035_o_0;
 wire n_10034_o_0;
 wire n_10033_o_0;
 wire n_10032_o_0;
 wire n_10031_o_0;
 wire n_10030_o_0;
 wire n_10029_o_0;
 wire n_10028_o_0;
 wire n_10027_o_0;
 wire n_10026_o_0;
 wire n_10025_o_0;
 wire n_10024_o_0;
 wire n_10023_o_0;
 wire n_10022_o_0;
 wire n_10021_o_0;
 wire n_10020_o_0;
 wire n_10019_o_0;
 wire n_10018_o_0;
 wire n_10017_o_0;
 wire n_10016_o_0;
 wire n_10015_o_0;
 wire n_10014_o_0;
 wire n_10013_o_0;
 wire n_10012_o_0;
 wire n_10011_o_0;
 wire n_10010_o_0;
 wire n_10009_o_0;
 wire n_10008_o_0;
 wire n_10007_o_0;
 wire n_10006_o_0;
 wire n_10005_o_0;
 wire n_10004_o_0;
 wire n_10003_o_0;
 wire n_10002_o_0;
 wire n_10001_o_0;
 wire n_10000_o_0;
 wire n_9999_o_0;
 wire n_9998_o_0;
 wire n_9997_o_0;
 wire n_9996_o_0;
 wire n_9995_o_0;
 wire n_9994_o_0;
 wire n_9993_o_0;
 wire n_9992_o_0;
 wire n_9991_o_0;
 wire n_9990_o_0;
 wire n_9989_o_0;
 wire n_9988_o_0;
 wire n_9987_o_0;
 wire n_9986_o_0;
 wire n_9985_o_0;
 wire n_9984_o_0;
 wire n_9983_o_0;
 wire n_9982_o_0;
 wire n_9981_o_0;
 wire n_9980_o_0;
 wire n_9979_o_0;
 wire n_9978_o_0;
 wire n_9977_o_0;
 wire n_9976_o_0;
 wire n_9975_o_0;
 wire n_9974_o_0;
 wire n_9973_o_0;
 wire n_9972_o_0;
 wire n_9971_o_0;
 wire n_9970_o_0;
 wire n_9969_o_0;
 wire n_9968_o_0;
 wire n_9967_o_0;
 wire n_9966_o_0;
 wire n_9965_o_0;
 wire n_9964_o_0;
 wire n_9963_o_0;
 wire n_9962_o_0;
 wire n_9961_o_0;
 wire n_9960_o_0;
 wire n_9959_o_0;
 wire n_9958_o_0;
 wire n_9957_o_0;
 wire n_9956_o_0;
 wire n_9955_o_0;
 wire n_9954_o_0;
 wire n_9953_o_0;
 wire n_9952_o_0;
 wire n_9951_o_0;
 wire n_9950_o_0;
 wire n_9949_o_0;
 wire n_9948_o_0;
 wire n_9947_o_0;
 wire n_9946_o_0;
 wire n_9945_o_0;
 wire n_9944_o_0;
 wire n_9943_o_0;
 wire n_9942_o_0;
 wire n_9941_o_0;
 wire n_9940_o_0;
 wire n_9939_o_0;
 wire n_9938_o_0;
 wire n_9937_o_0;
 wire n_9936_o_0;
 wire n_9935_o_0;
 wire n_9934_o_0;
 wire n_9933_o_0;
 wire n_9932_o_0;
 wire n_9931_o_0;
 wire n_9930_o_0;
 wire n_9929_o_0;
 wire n_9928_o_0;
 wire n_9927_o_0;
 wire n_9926_o_0;
 wire n_9925_o_0;
 wire n_9924_o_0;
 wire n_9923_o_0;
 wire n_9922_o_0;
 wire n_9921_o_0;
 wire n_9920_o_0;
 wire n_9919_o_0;
 wire n_9918_o_0;
 wire n_9917_o_0;
 wire n_9916_o_0;
 wire n_9915_o_0;
 wire n_9914_o_0;
 wire n_9913_o_0;
 wire n_9912_o_0;
 wire n_9911_o_0;
 wire n_9910_o_0;
 wire n_9909_o_0;
 wire n_9908_o_0;
 wire n_9907_o_0;
 wire n_9906_o_0;
 wire n_9905_o_0;
 wire n_9904_o_0;
 wire n_9903_o_0;
 wire n_9902_o_0;
 wire n_9901_o_0;
 wire n_9900_o_0;
 wire n_9899_o_0;
 wire n_9898_o_0;
 wire n_9897_o_0;
 wire n_9896_o_0;
 wire n_9895_o_0;
 wire n_9894_o_0;
 wire n_9893_o_0;
 wire n_9892_o_0;
 wire n_9891_o_0;
 wire n_9890_o_0;
 wire n_9889_o_0;
 wire n_9888_o_0;
 wire n_9887_o_0;
 wire n_9886_o_0;
 wire n_9885_o_0;
 wire n_9884_o_0;
 wire n_9883_o_0;
 wire n_9882_o_0;
 wire n_9881_o_0;
 wire n_9880_o_0;
 wire n_9879_o_0;
 wire n_9878_o_0;
 wire n_9877_o_0;
 wire n_9876_o_0;
 wire n_9875_o_0;
 wire n_9874_o_0;
 wire n_9873_o_0;
 wire n_9872_o_0;
 wire n_9871_o_0;
 wire n_9870_o_0;
 wire n_9869_o_0;
 wire n_9868_o_0;
 wire n_9867_o_0;
 wire n_9866_o_0;
 wire n_9865_o_0;
 wire n_9864_o_0;
 wire n_9863_o_0;
 wire n_9862_o_0;
 wire n_9861_o_0;
 wire n_9860_o_0;
 wire n_9859_o_0;
 wire n_9858_o_0;
 wire n_9857_o_0;
 wire n_9856_o_0;
 wire n_9855_o_0;
 wire n_9854_o_0;
 wire n_9853_o_0;
 wire n_9852_o_0;
 wire n_9851_o_0;
 wire n_9850_o_0;
 wire n_9849_o_0;
 wire n_9848_o_0;
 wire n_9847_o_0;
 wire n_9846_o_0;
 wire n_9845_o_0;
 wire n_9844_o_0;
 wire n_9843_o_0;
 wire n_9842_o_0;
 wire n_9841_o_0;
 wire n_9840_o_0;
 wire n_9839_o_0;
 wire n_9838_o_0;
 wire n_9837_o_0;
 wire n_9836_o_0;
 wire n_9835_o_0;
 wire n_9834_o_0;
 wire n_9833_o_0;
 wire n_9832_o_0;
 wire n_9831_o_0;
 wire n_9830_o_0;
 wire n_9829_o_0;
 wire n_9828_o_0;
 wire n_9827_o_0;
 wire n_9826_o_0;
 wire n_9825_o_0;
 wire n_9824_o_0;
 wire n_9823_o_0;
 wire n_9822_o_0;
 wire n_9821_o_0;
 wire n_9820_o_0;
 wire n_9819_o_0;
 wire n_9818_o_0;
 wire n_9817_o_0;
 wire n_9816_o_0;
 wire n_9815_o_0;
 wire n_9814_o_0;
 wire n_9813_o_0;
 wire n_9812_o_0;
 wire n_9811_o_0;
 wire n_9810_o_0;
 wire n_9809_o_0;
 wire n_9808_o_0;
 wire n_9807_o_0;
 wire n_9806_o_0;
 wire n_9805_o_0;
 wire n_9804_o_0;
 wire n_9803_o_0;
 wire n_9802_o_0;
 wire n_9801_o_0;
 wire n_9800_o_0;
 wire n_9799_o_0;
 wire n_9798_o_0;
 wire n_9797_o_0;
 wire n_9796_o_0;
 wire n_9795_o_0;
 wire n_9794_o_0;
 wire n_9793_o_0;
 wire n_9792_o_0;
 wire n_9791_o_0;
 wire n_9790_o_0;
 wire n_9789_o_0;
 wire n_9788_o_0;
 wire n_9787_o_0;
 wire n_9786_o_0;
 wire n_9785_o_0;
 wire n_9784_o_0;
 wire n_9783_o_0;
 wire n_9782_o_0;
 wire n_9781_o_0;
 wire n_9780_o_0;
 wire n_9779_o_0;
 wire n_9778_o_0;
 wire n_9777_o_0;
 wire n_9776_o_0;
 wire n_9775_o_0;
 wire n_9774_o_0;
 wire n_9773_o_0;
 wire n_9772_o_0;
 wire n_9771_o_0;
 wire n_9770_o_0;
 wire n_9769_o_0;
 wire n_9768_o_0;
 wire n_9767_o_0;
 wire n_9766_o_0;
 wire n_9765_o_0;
 wire n_9764_o_0;
 wire n_9763_o_0;
 wire n_9762_o_0;
 wire n_9761_o_0;
 wire n_9760_o_0;
 wire n_9759_o_0;
 wire n_9758_o_0;
 wire n_9757_o_0;
 wire n_9756_o_0;
 wire n_9755_o_0;
 wire n_9754_o_0;
 wire n_9753_o_0;
 wire n_9752_o_0;
 wire n_9751_o_0;
 wire n_9750_o_0;
 wire n_9749_o_0;
 wire n_9748_o_0;
 wire n_9747_o_0;
 wire n_9746_o_0;
 wire n_9745_o_0;
 wire n_9744_o_0;
 wire n_9743_o_0;
 wire n_9742_o_0;
 wire n_9741_o_0;
 wire n_9740_o_0;
 wire n_9739_o_0;
 wire n_9738_o_0;
 wire n_9737_o_0;
 wire n_9736_o_0;
 wire n_9735_o_0;
 wire n_9734_o_0;
 wire n_9733_o_0;
 wire n_9732_o_0;
 wire n_9731_o_0;
 wire n_9730_o_0;
 wire n_9729_o_0;
 wire n_9728_o_0;
 wire n_9727_o_0;
 wire n_9726_o_0;
 wire n_9725_o_0;
 wire n_9724_o_0;
 wire n_9723_o_0;
 wire n_9722_o_0;
 wire n_9721_o_0;
 wire n_9720_o_0;
 wire n_9719_o_0;
 wire n_9718_o_0;
 wire n_9717_o_0;
 wire n_9716_o_0;
 wire n_9715_o_0;
 wire n_9714_o_0;
 wire n_9713_o_0;
 wire n_9712_o_0;
 wire n_9711_o_0;
 wire n_9710_o_0;
 wire n_9709_o_0;
 wire n_9708_o_0;
 wire n_9707_o_0;
 wire n_9706_o_0;
 wire n_9705_o_0;
 wire n_9704_o_0;
 wire n_9703_o_0;
 wire n_9702_o_0;
 wire n_9701_o_0;
 wire n_9700_o_0;
 wire n_9699_o_0;
 wire n_9698_o_0;
 wire n_9697_o_0;
 wire n_9696_o_0;
 wire n_9695_o_0;
 wire n_9694_o_0;
 wire n_9693_o_0;
 wire n_9692_o_0;
 wire n_9691_o_0;
 wire n_9690_o_0;
 wire n_9689_o_0;
 wire n_9688_o_0;
 wire n_9687_o_0;
 wire n_9686_o_0;
 wire n_9685_o_0;
 wire n_9684_o_0;
 wire n_9683_o_0;
 wire n_9682_o_0;
 wire n_9681_o_0;
 wire n_9680_o_0;
 wire n_9679_o_0;
 wire n_9678_o_0;
 wire n_9677_o_0;
 wire n_9676_o_0;
 wire n_9675_o_0;
 wire n_9674_o_0;
 wire n_9673_o_0;
 wire n_9672_o_0;
 wire n_9671_o_0;
 wire n_9670_o_0;
 wire n_9669_o_0;
 wire n_9668_o_0;
 wire n_9667_o_0;
 wire n_9666_o_0;
 wire n_9665_o_0;
 wire n_9664_o_0;
 wire n_9663_o_0;
 wire n_9662_o_0;
 wire n_9661_o_0;
 wire n_9660_o_0;
 wire n_9659_o_0;
 wire n_9658_o_0;
 wire n_9657_o_0;
 wire n_9656_o_0;
 wire n_9655_o_0;
 wire n_9654_o_0;
 wire n_9653_o_0;
 wire n_9652_o_0;
 wire n_9651_o_0;
 wire n_9650_o_0;
 wire n_9649_o_0;
 wire n_9648_o_0;
 wire n_9647_o_0;
 wire n_9646_o_0;
 wire n_9645_o_0;
 wire n_9644_o_0;
 wire n_9643_o_0;
 wire n_9642_o_0;
 wire n_9641_o_0;
 wire n_9640_o_0;
 wire n_9639_o_0;
 wire n_9638_o_0;
 wire n_9637_o_0;
 wire n_9636_o_0;
 wire n_9635_o_0;
 wire n_9634_o_0;
 wire n_9633_o_0;
 wire n_9632_o_0;
 wire n_9631_o_0;
 wire n_9630_o_0;
 wire n_9629_o_0;
 wire n_9628_o_0;
 wire n_9627_o_0;
 wire n_9626_o_0;
 wire n_9625_o_0;
 wire n_9624_o_0;
 wire n_9623_o_0;
 wire n_9622_o_0;
 wire n_9621_o_0;
 wire n_9620_o_0;
 wire n_9619_o_0;
 wire n_9618_o_0;
 wire n_9617_o_0;
 wire n_9616_o_0;
 wire n_9615_o_0;
 wire n_9614_o_0;
 wire n_9613_o_0;
 wire n_9612_o_0;
 wire n_9611_o_0;
 wire n_9610_o_0;
 wire n_9609_o_0;
 wire n_9608_o_0;
 wire n_9607_o_0;
 wire n_9606_o_0;
 wire n_9605_o_0;
 wire n_9604_o_0;
 wire n_9603_o_0;
 wire n_9602_o_0;
 wire n_9601_o_0;
 wire n_9600_o_0;
 wire n_9599_o_0;
 wire n_9598_o_0;
 wire n_9597_o_0;
 wire n_9596_o_0;
 wire n_9595_o_0;
 wire n_9594_o_0;
 wire n_9593_o_0;
 wire n_9592_o_0;
 wire n_9591_o_0;
 wire n_9590_o_0;
 wire n_9589_o_0;
 wire n_9588_o_0;
 wire n_9587_o_0;
 wire n_9586_o_0;
 wire n_9585_o_0;
 wire n_9584_o_0;
 wire n_9583_o_0;
 wire n_9582_o_0;
 wire n_9581_o_0;
 wire n_9580_o_0;
 wire n_9579_o_0;
 wire n_9578_o_0;
 wire n_9577_o_0;
 wire n_9576_o_0;
 wire n_9575_o_0;
 wire n_9574_o_0;
 wire n_9573_o_0;
 wire n_9572_o_0;
 wire n_9571_o_0;
 wire n_9570_o_0;
 wire n_9569_o_0;
 wire n_9568_o_0;
 wire n_9567_o_0;
 wire n_9566_o_0;
 wire n_9565_o_0;
 wire n_9564_o_0;
 wire n_9563_o_0;
 wire n_9562_o_0;
 wire n_9561_o_0;
 wire n_9560_o_0;
 wire n_9559_o_0;
 wire n_9558_o_0;
 wire n_9557_o_0;
 wire n_9556_o_0;
 wire n_9555_o_0;
 wire n_9554_o_0;
 wire n_9553_o_0;
 wire n_9552_o_0;
 wire n_9551_o_0;
 wire n_9550_o_0;
 wire n_9549_o_0;
 wire n_9548_o_0;
 wire n_9547_o_0;
 wire n_9546_o_0;
 wire n_9545_o_0;
 wire n_9544_o_0;
 wire n_9543_o_0;
 wire n_9542_o_0;
 wire n_9541_o_0;
 wire n_9540_o_0;
 wire n_9539_o_0;
 wire n_9538_o_0;
 wire n_9537_o_0;
 wire n_9536_o_0;
 wire n_9535_o_0;
 wire n_9534_o_0;
 wire n_9533_o_0;
 wire n_9532_o_0;
 wire n_9531_o_0;
 wire n_9530_o_0;
 wire n_9529_o_0;
 wire n_9528_o_0;
 wire n_9527_o_0;
 wire n_9526_o_0;
 wire n_9525_o_0;
 wire n_9524_o_0;
 wire n_9523_o_0;
 wire n_9522_o_0;
 wire n_9521_o_0;
 wire n_9520_o_0;
 wire n_9519_o_0;
 wire n_9518_o_0;
 wire n_9517_o_0;
 wire n_9516_o_0;
 wire n_9515_o_0;
 wire n_9514_o_0;
 wire n_9513_o_0;
 wire n_9512_o_0;
 wire n_9511_o_0;
 wire n_9510_o_0;
 wire n_9509_o_0;
 wire n_9508_o_0;
 wire n_9507_o_0;
 wire n_9506_o_0;
 wire n_9505_o_0;
 wire n_9504_o_0;
 wire n_9503_o_0;
 wire n_9502_o_0;
 wire n_9501_o_0;
 wire n_9500_o_0;
 wire n_9499_o_0;
 wire n_9498_o_0;
 wire n_9497_o_0;
 wire n_9496_o_0;
 wire n_9495_o_0;
 wire n_9494_o_0;
 wire n_9493_o_0;
 wire n_9492_o_0;
 wire n_9491_o_0;
 wire n_9490_o_0;
 wire n_9489_o_0;
 wire n_9488_o_0;
 wire n_9487_o_0;
 wire n_9486_o_0;
 wire n_9485_o_0;
 wire n_9484_o_0;
 wire n_9483_o_0;
 wire n_9482_o_0;
 wire n_9481_o_0;
 wire n_9480_o_0;
 wire n_9479_o_0;
 wire n_9478_o_0;
 wire n_9477_o_0;
 wire n_9476_o_0;
 wire n_9475_o_0;
 wire n_9474_o_0;
 wire n_9473_o_0;
 wire n_9472_o_0;
 wire n_9471_o_0;
 wire n_9470_o_0;
 wire n_9469_o_0;
 wire n_9468_o_0;
 wire n_9467_o_0;
 wire n_9466_o_0;
 wire n_9465_o_0;
 wire n_9464_o_0;
 wire n_9463_o_0;
 wire n_9462_o_0;
 wire n_9461_o_0;
 wire n_9460_o_0;
 wire n_9459_o_0;
 wire n_9458_o_0;
 wire n_9457_o_0;
 wire n_9456_o_0;
 wire n_9455_o_0;
 wire n_9454_o_0;
 wire n_9453_o_0;
 wire n_9452_o_0;
 wire n_9451_o_0;
 wire n_9450_o_0;
 wire n_9449_o_0;
 wire n_9448_o_0;
 wire n_9447_o_0;
 wire n_9446_o_0;
 wire n_9445_o_0;
 wire n_9444_o_0;
 wire n_9443_o_0;
 wire n_9442_o_0;
 wire n_9441_o_0;
 wire n_9440_o_0;
 wire n_9439_o_0;
 wire n_9438_o_0;
 wire n_9437_o_0;
 wire n_9436_o_0;
 wire n_9435_o_0;
 wire n_9434_o_0;
 wire n_9433_o_0;
 wire n_9432_o_0;
 wire n_9431_o_0;
 wire n_9430_o_0;
 wire n_9429_o_0;
 wire n_9428_o_0;
 wire n_9427_o_0;
 wire n_9426_o_0;
 wire n_9425_o_0;
 wire n_9424_o_0;
 wire n_9423_o_0;
 wire n_9422_o_0;
 wire n_9421_o_0;
 wire n_9420_o_0;
 wire n_9419_o_0;
 wire n_9418_o_0;
 wire n_9417_o_0;
 wire n_9416_o_1;
 wire n_9416_o_0;
 wire n_9415_o_0;
 wire n_9414_o_0;
 wire n_9413_o_0;
 wire n_9412_o_0;
 wire n_9411_o_0;
 wire n_9410_o_0;
 wire n_9409_o_0;
 wire n_9408_o_0;
 wire n_9407_o_0;
 wire n_9406_o_0;
 wire n_9405_o_0;
 wire n_9404_o_0;
 wire n_9403_o_0;
 wire n_9402_o_0;
 wire n_9401_o_0;
 wire n_9400_o_0;
 wire n_9399_o_0;
 wire n_9398_o_0;
 wire n_9397_o_0;
 wire n_9396_o_0;
 wire n_9395_o_0;
 wire n_9394_o_0;
 wire n_9393_o_0;
 wire n_9392_o_0;
 wire n_9391_o_0;
 wire n_9390_o_0;
 wire n_9389_o_0;
 wire n_9388_o_0;
 wire n_9387_o_0;
 wire n_9386_o_0;
 wire n_9385_o_0;
 wire n_9384_o_0;
 wire n_9383_o_0;
 wire n_9382_o_0;
 wire n_9381_o_0;
 wire n_9380_o_0;
 wire n_9379_o_0;
 wire n_9378_o_0;
 wire n_9377_o_0;
 wire n_9376_o_0;
 wire n_9375_o_0;
 wire n_9374_o_0;
 wire n_9373_o_0;
 wire n_9372_o_0;
 wire n_9371_o_0;
 wire n_9370_o_0;
 wire n_9369_o_0;
 wire n_9368_o_0;
 wire n_9367_o_0;
 wire n_9366_o_0;
 wire n_9365_o_0;
 wire n_9364_o_0;
 wire n_9363_o_0;
 wire n_9362_o_0;
 wire n_9361_o_0;
 wire n_9360_o_0;
 wire n_9359_o_0;
 wire n_9358_o_0;
 wire n_9357_o_0;
 wire n_9356_o_0;
 wire n_9355_o_0;
 wire n_9354_o_0;
 wire n_9353_o_0;
 wire n_9352_o_0;
 wire n_9351_o_0;
 wire n_9350_o_0;
 wire n_9349_o_0;
 wire n_9348_o_0;
 wire n_9347_o_0;
 wire n_9346_o_0;
 wire n_9345_o_0;
 wire n_9344_o_0;
 wire n_9343_o_0;
 wire n_9342_o_0;
 wire n_9341_o_0;
 wire n_9340_o_0;
 wire n_9339_o_0;
 wire n_9338_o_0;
 wire n_9337_o_0;
 wire n_9336_o_0;
 wire n_9335_o_0;
 wire n_9334_o_0;
 wire n_9333_o_0;
 wire n_9332_o_0;
 wire n_9331_o_0;
 wire n_9330_o_0;
 wire n_9329_o_0;
 wire n_9328_o_0;
 wire n_9327_o_0;
 wire n_9326_o_0;
 wire n_9325_o_0;
 wire n_9324_o_0;
 wire n_9323_o_0;
 wire n_9322_o_0;
 wire n_9321_o_0;
 wire n_9320_o_0;
 wire n_9319_o_0;
 wire n_9318_o_0;
 wire n_9317_o_0;
 wire n_9316_o_0;
 wire n_9315_o_0;
 wire n_9314_o_0;
 wire n_9313_o_0;
 wire n_9312_o_0;
 wire n_9311_o_0;
 wire n_9310_o_0;
 wire n_9309_o_0;
 wire n_9308_o_0;
 wire n_9307_o_0;
 wire n_9306_o_0;
 wire n_9305_o_0;
 wire n_9304_o_0;
 wire n_9303_o_0;
 wire n_9302_o_0;
 wire n_9301_o_0;
 wire n_9300_o_0;
 wire n_9299_o_0;
 wire n_9298_o_0;
 wire n_9297_o_0;
 wire n_9296_o_0;
 wire n_9295_o_0;
 wire n_9294_o_0;
 wire n_9293_o_0;
 wire n_9292_o_0;
 wire n_9291_o_0;
 wire n_9290_o_0;
 wire n_9289_o_0;
 wire n_9288_o_0;
 wire n_9287_o_0;
 wire n_9286_o_0;
 wire n_9285_o_0;
 wire n_9284_o_0;
 wire n_9283_o_0;
 wire n_9282_o_0;
 wire n_9281_o_0;
 wire n_9280_o_0;
 wire n_9279_o_0;
 wire n_9278_o_0;
 wire n_9277_o_0;
 wire n_9276_o_0;
 wire n_9275_o_0;
 wire n_9274_o_0;
 wire n_9273_o_0;
 wire n_9272_o_0;
 wire n_9271_o_0;
 wire n_9270_o_0;
 wire n_9269_o_0;
 wire n_9268_o_0;
 wire n_9267_o_0;
 wire n_9266_o_0;
 wire n_9265_o_0;
 wire n_9264_o_0;
 wire n_9263_o_0;
 wire n_9262_o_0;
 wire n_9261_o_0;
 wire n_9260_o_0;
 wire n_9259_o_0;
 wire n_9258_o_0;
 wire n_9257_o_0;
 wire n_9256_o_0;
 wire n_9255_o_0;
 wire n_9254_o_0;
 wire n_9253_o_0;
 wire n_9252_o_0;
 wire n_9251_o_0;
 wire n_9250_o_0;
 wire n_9249_o_0;
 wire n_9248_o_0;
 wire n_9247_o_0;
 wire n_9246_o_0;
 wire n_9245_o_0;
 wire n_9244_o_0;
 wire n_9243_o_0;
 wire n_9242_o_0;
 wire n_9241_o_0;
 wire n_9240_o_0;
 wire n_9239_o_0;
 wire n_9238_o_0;
 wire n_9237_o_0;
 wire n_9236_o_0;
 wire n_9235_o_0;
 wire n_9234_o_0;
 wire n_9233_o_0;
 wire n_9232_o_0;
 wire n_9231_o_0;
 wire n_9230_o_0;
 wire n_9229_o_0;
 wire n_9228_o_0;
 wire n_9227_o_0;
 wire n_9226_o_0;
 wire n_9225_o_0;
 wire n_9224_o_0;
 wire n_9223_o_0;
 wire n_9222_o_0;
 wire n_9221_o_0;
 wire n_9220_o_0;
 wire n_9219_o_0;
 wire n_9218_o_0;
 wire n_9217_o_0;
 wire n_9216_o_0;
 wire n_9215_o_0;
 wire n_9214_o_0;
 wire n_9213_o_0;
 wire n_9212_o_0;
 wire n_9211_o_0;
 wire n_9210_o_0;
 wire n_9209_o_0;
 wire n_9208_o_0;
 wire n_9207_o_0;
 wire n_9206_o_0;
 wire n_9205_o_0;
 wire n_9204_o_0;
 wire n_9203_o_0;
 wire n_9202_o_0;
 wire n_9201_o_0;
 wire n_9200_o_0;
 wire n_9199_o_0;
 wire n_9198_o_0;
 wire n_9197_o_0;
 wire n_9196_o_0;
 wire n_9195_o_0;
 wire n_9194_o_0;
 wire n_9193_o_0;
 wire n_9192_o_0;
 wire n_9191_o_0;
 wire n_9190_o_0;
 wire n_9189_o_0;
 wire n_9188_o_0;
 wire n_9187_o_0;
 wire n_9186_o_0;
 wire n_9185_o_0;
 wire n_9184_o_0;
 wire n_9183_o_0;
 wire n_9182_o_0;
 wire n_9181_o_0;
 wire n_9180_o_0;
 wire n_9179_o_0;
 wire n_9178_o_0;
 wire n_9177_o_0;
 wire n_9176_o_0;
 wire n_9175_o_0;
 wire n_9174_o_0;
 wire n_9173_o_0;
 wire n_9172_o_0;
 wire n_9171_o_0;
 wire n_9170_o_0;
 wire n_9169_o_0;
 wire n_9168_o_0;
 wire n_9167_o_0;
 wire n_9166_o_0;
 wire n_9165_o_0;
 wire n_9164_o_0;
 wire n_9163_o_0;
 wire n_9162_o_0;
 wire n_9161_o_0;
 wire n_9160_o_0;
 wire n_9159_o_0;
 wire n_9158_o_0;
 wire n_9157_o_0;
 wire n_9156_o_0;
 wire n_9155_o_0;
 wire n_9154_o_0;
 wire n_9153_o_0;
 wire n_9152_o_0;
 wire n_9151_o_0;
 wire n_9150_o_0;
 wire n_9149_o_0;
 wire n_9148_o_0;
 wire n_9147_o_0;
 wire n_9146_o_0;
 wire n_9145_o_0;
 wire n_9144_o_0;
 wire n_9143_o_0;
 wire n_9142_o_0;
 wire n_9141_o_0;
 wire n_9140_o_0;
 wire n_9139_o_0;
 wire n_9138_o_0;
 wire n_9137_o_0;
 wire n_9136_o_0;
 wire n_9135_o_0;
 wire n_9134_o_0;
 wire n_9133_o_0;
 wire n_9132_o_0;
 wire n_9131_o_0;
 wire n_9130_o_0;
 wire n_9129_o_0;
 wire n_9128_o_0;
 wire n_9127_o_0;
 wire n_9126_o_0;
 wire n_9125_o_0;
 wire n_9124_o_0;
 wire n_9123_o_0;
 wire n_9122_o_0;
 wire n_9121_o_0;
 wire n_9120_o_0;
 wire n_9119_o_0;
 wire n_9118_o_0;
 wire n_9117_o_0;
 wire n_9116_o_0;
 wire n_9115_o_0;
 wire n_9114_o_0;
 wire n_9113_o_0;
 wire n_9112_o_0;
 wire n_9111_o_0;
 wire n_9110_o_0;
 wire n_9109_o_0;
 wire n_9108_o_0;
 wire n_9107_o_0;
 wire n_9106_o_0;
 wire n_9105_o_0;
 wire n_9104_o_0;
 wire n_9103_o_0;
 wire n_9102_o_0;
 wire n_9101_o_0;
 wire n_9100_o_0;
 wire n_9099_o_0;
 wire n_9098_o_0;
 wire n_9097_o_0;
 wire n_9096_o_0;
 wire n_9095_o_0;
 wire n_9094_o_0;
 wire n_9093_o_0;
 wire n_9092_o_0;
 wire n_9091_o_0;
 wire n_9090_o_0;
 wire n_9089_o_0;
 wire n_9088_o_0;
 wire n_9087_o_0;
 wire n_9086_o_0;
 wire n_9085_o_0;
 wire n_9084_o_0;
 wire n_9083_o_0;
 wire n_9082_o_0;
 wire n_9081_o_0;
 wire n_9080_o_0;
 wire n_9079_o_0;
 wire n_9078_o_0;
 wire n_9077_o_0;
 wire n_9076_o_0;
 wire n_9075_o_0;
 wire n_9074_o_0;
 wire n_9073_o_0;
 wire n_9072_o_0;
 wire n_9071_o_0;
 wire n_9070_o_0;
 wire n_9069_o_0;
 wire n_9068_o_0;
 wire n_9067_o_0;
 wire n_9066_o_0;
 wire n_9065_o_0;
 wire n_9064_o_0;
 wire n_9063_o_0;
 wire n_9062_o_0;
 wire n_9061_o_0;
 wire n_9060_o_0;
 wire n_9059_o_0;
 wire n_9058_o_0;
 wire n_9057_o_0;
 wire n_9056_o_0;
 wire n_9055_o_0;
 wire n_9054_o_0;
 wire n_9053_o_0;
 wire n_9052_o_0;
 wire n_9051_o_0;
 wire n_9050_o_0;
 wire n_9049_o_0;
 wire n_9048_o_0;
 wire n_9047_o_0;
 wire n_9046_o_0;
 wire n_9045_o_0;
 wire n_9044_o_0;
 wire n_9043_o_0;
 wire n_9042_o_0;
 wire n_9041_o_0;
 wire n_9040_o_0;
 wire n_9039_o_0;
 wire n_9038_o_0;
 wire n_9037_o_0;
 wire n_9036_o_0;
 wire n_9035_o_0;
 wire n_9034_o_0;
 wire n_9033_o_0;
 wire n_9032_o_0;
 wire n_9031_o_0;
 wire n_9030_o_0;
 wire n_9029_o_0;
 wire n_9028_o_0;
 wire n_9027_o_0;
 wire n_9026_o_0;
 wire n_9025_o_0;
 wire n_9024_o_0;
 wire n_9023_o_0;
 wire n_9022_o_0;
 wire n_9021_o_0;
 wire n_9020_o_0;
 wire n_9019_o_0;
 wire n_9018_o_0;
 wire n_9017_o_0;
 wire n_9016_o_0;
 wire n_9015_o_0;
 wire n_9014_o_0;
 wire n_9013_o_0;
 wire n_9012_o_0;
 wire n_9011_o_0;
 wire n_9010_o_0;
 wire n_9009_o_0;
 wire n_9008_o_0;
 wire n_9007_o_0;
 wire n_9006_o_0;
 wire n_9005_o_0;
 wire n_9004_o_0;
 wire n_9003_o_0;
 wire n_9002_o_0;
 wire n_9001_o_0;
 wire n_9000_o_0;
 wire n_8999_o_0;
 wire n_8998_o_0;
 wire n_8997_o_0;
 wire n_8996_o_0;
 wire n_8995_o_0;
 wire n_8994_o_0;
 wire n_8993_o_0;
 wire n_8992_o_0;
 wire n_8991_o_0;
 wire n_8990_o_0;
 wire n_8989_o_0;
 wire n_8988_o_0;
 wire n_8987_o_0;
 wire n_8986_o_0;
 wire n_8985_o_0;
 wire n_8984_o_0;
 wire n_8983_o_0;
 wire n_8982_o_0;
 wire n_8981_o_0;
 wire n_8980_o_0;
 wire n_8979_o_0;
 wire n_8978_o_0;
 wire n_8977_o_0;
 wire n_8976_o_0;
 wire n_8975_o_0;
 wire n_8974_o_0;
 wire n_8973_o_0;
 wire n_8972_o_0;
 wire n_8971_o_0;
 wire n_8970_o_0;
 wire n_8969_o_0;
 wire n_8968_o_0;
 wire n_8967_o_0;
 wire n_8966_o_0;
 wire n_8965_o_0;
 wire n_8964_o_0;
 wire n_8963_o_0;
 wire n_8962_o_0;
 wire n_8961_o_0;
 wire n_8960_o_0;
 wire n_8959_o_0;
 wire n_8958_o_0;
 wire n_8957_o_0;
 wire n_8956_o_0;
 wire n_8955_o_0;
 wire n_8954_o_0;
 wire n_8953_o_0;
 wire n_8952_o_0;
 wire n_8951_o_0;
 wire n_8950_o_0;
 wire n_8949_o_0;
 wire n_8948_o_0;
 wire n_8947_o_0;
 wire n_8946_o_0;
 wire n_8945_o_0;
 wire n_8944_o_0;
 wire n_8943_o_0;
 wire n_8942_o_0;
 wire n_8941_o_0;
 wire n_8940_o_0;
 wire n_8939_o_0;
 wire n_8938_o_0;
 wire n_8937_o_0;
 wire n_8936_o_0;
 wire n_8935_o_0;
 wire n_8934_o_0;
 wire n_8933_o_0;
 wire n_8932_o_0;
 wire n_8931_o_0;
 wire n_8930_o_0;
 wire n_8929_o_0;
 wire n_8928_o_0;
 wire n_8927_o_0;
 wire n_8926_o_0;
 wire n_8925_o_0;
 wire n_8924_o_0;
 wire n_8923_o_0;
 wire n_8922_o_0;
 wire n_8921_o_0;
 wire n_8920_o_0;
 wire n_8919_o_0;
 wire n_8918_o_0;
 wire n_8917_o_0;
 wire n_8916_o_0;
 wire n_8915_o_0;
 wire n_8914_o_0;
 wire n_8913_o_0;
 wire n_8912_o_0;
 wire n_8911_o_0;
 wire n_8910_o_0;
 wire n_8909_o_0;
 wire n_8908_o_0;
 wire n_8907_o_0;
 wire n_8906_o_0;
 wire n_8905_o_0;
 wire n_8904_o_0;
 wire n_8903_o_0;
 wire n_8902_o_0;
 wire n_8901_o_0;
 wire n_8900_o_0;
 wire n_8899_o_0;
 wire n_8898_o_0;
 wire n_8897_o_0;
 wire n_8896_o_0;
 wire n_8895_o_0;
 wire n_8894_o_0;
 wire n_8893_o_0;
 wire n_8892_o_0;
 wire n_8891_o_0;
 wire n_8890_o_0;
 wire n_8889_o_0;
 wire n_8888_o_0;
 wire n_8887_o_0;
 wire n_8886_o_0;
 wire n_8885_o_0;
 wire n_8884_o_0;
 wire n_8883_o_0;
 wire n_8882_o_0;
 wire n_8881_o_0;
 wire n_8880_o_0;
 wire n_8879_o_0;
 wire n_8878_o_0;
 wire n_8877_o_0;
 wire n_8876_o_0;
 wire n_8875_o_0;
 wire n_8874_o_0;
 wire n_8873_o_0;
 wire n_8872_o_0;
 wire n_8871_o_0;
 wire n_8870_o_0;
 wire n_8869_o_0;
 wire n_8868_o_0;
 wire n_8867_o_0;
 wire n_8866_o_0;
 wire n_8865_o_0;
 wire n_8864_o_0;
 wire n_8863_o_0;
 wire n_8862_o_0;
 wire n_8861_o_0;
 wire n_8860_o_0;
 wire n_8859_o_0;
 wire n_8858_o_0;
 wire n_8857_o_0;
 wire n_8856_o_0;
 wire n_8855_o_0;
 wire n_8854_o_0;
 wire n_8853_o_0;
 wire n_8852_o_0;
 wire n_8851_o_0;
 wire n_8850_o_0;
 wire n_8849_o_0;
 wire n_8848_o_0;
 wire n_8847_o_0;
 wire n_8846_o_0;
 wire n_8845_o_0;
 wire n_8844_o_0;
 wire n_8843_o_0;
 wire n_8842_o_0;
 wire n_8841_o_0;
 wire n_8840_o_0;
 wire n_8839_o_0;
 wire n_8838_o_0;
 wire n_8837_o_0;
 wire n_8836_o_0;
 wire n_8835_o_0;
 wire n_8834_o_0;
 wire n_8833_o_0;
 wire n_8832_o_0;
 wire n_8831_o_0;
 wire n_8830_o_0;
 wire n_8829_o_0;
 wire n_8828_o_0;
 wire n_8827_o_0;
 wire n_8826_o_0;
 wire n_8825_o_0;
 wire n_8824_o_0;
 wire n_8823_o_0;
 wire n_8822_o_0;
 wire n_8821_o_0;
 wire n_8820_o_0;
 wire n_8819_o_0;
 wire n_8818_o_0;
 wire n_8817_o_0;
 wire n_8816_o_0;
 wire n_8815_o_0;
 wire n_8814_o_0;
 wire n_8813_o_0;
 wire n_8812_o_0;
 wire n_8811_o_0;
 wire n_8810_o_0;
 wire n_8809_o_0;
 wire n_8808_o_0;
 wire n_8807_o_0;
 wire n_8806_o_0;
 wire n_8805_o_0;
 wire n_8804_o_0;
 wire n_8803_o_0;
 wire n_8802_o_0;
 wire n_8801_o_0;
 wire n_8800_o_0;
 wire n_8799_o_0;
 wire n_8798_o_0;
 wire n_8797_o_0;
 wire n_8796_o_0;
 wire n_8795_o_0;
 wire n_8794_o_0;
 wire n_8793_o_0;
 wire n_8792_o_0;
 wire n_8791_o_0;
 wire n_8790_o_0;
 wire n_8789_o_0;
 wire n_8788_o_0;
 wire n_8787_o_0;
 wire n_8786_o_0;
 wire n_8785_o_0;
 wire n_8784_o_0;
 wire n_8783_o_0;
 wire n_8782_o_0;
 wire n_8781_o_0;
 wire n_8780_o_0;
 wire n_8779_o_0;
 wire n_8778_o_0;
 wire n_8777_o_0;
 wire n_8776_o_0;
 wire n_8775_o_0;
 wire n_8774_o_0;
 wire n_8773_o_0;
 wire n_8772_o_0;
 wire n_8771_o_0;
 wire n_8770_o_0;
 wire n_8769_o_0;
 wire n_8768_o_0;
 wire n_8767_o_0;
 wire n_8766_o_0;
 wire n_8765_o_0;
 wire n_8764_o_0;
 wire n_8763_o_0;
 wire n_8762_o_0;
 wire n_8761_o_0;
 wire n_8760_o_0;
 wire n_8759_o_0;
 wire n_8758_o_0;
 wire n_8757_o_0;
 wire n_8756_o_0;
 wire n_8755_o_0;
 wire n_8754_o_0;
 wire n_8753_o_0;
 wire n_8752_o_0;
 wire n_8751_o_0;
 wire n_8750_o_0;
 wire n_8749_o_0;
 wire n_8748_o_0;
 wire n_8747_o_0;
 wire n_8746_o_0;
 wire n_8745_o_0;
 wire n_8744_o_0;
 wire n_8743_o_0;
 wire n_8742_o_0;
 wire n_8741_o_0;
 wire n_8740_o_0;
 wire n_8739_o_0;
 wire n_8738_o_0;
 wire n_8737_o_0;
 wire n_8736_o_0;
 wire n_8735_o_0;
 wire n_8734_o_0;
 wire n_8733_o_0;
 wire n_8732_o_0;
 wire n_8731_o_0;
 wire n_8730_o_0;
 wire n_8729_o_0;
 wire n_8728_o_0;
 wire n_8727_o_0;
 wire n_8726_o_0;
 wire n_8725_o_0;
 wire n_8724_o_0;
 wire n_8723_o_0;
 wire n_8722_o_0;
 wire n_8721_o_0;
 wire n_8720_o_0;
 wire n_8719_o_0;
 wire n_8718_o_0;
 wire n_8717_o_0;
 wire n_8716_o_0;
 wire n_8715_o_0;
 wire n_8714_o_0;
 wire n_8713_o_0;
 wire n_8712_o_0;
 wire n_8711_o_0;
 wire n_8710_o_0;
 wire n_8709_o_0;
 wire n_8708_o_0;
 wire n_8707_o_0;
 wire n_8706_o_0;
 wire n_8705_o_0;
 wire n_8704_o_0;
 wire n_8703_o_0;
 wire n_8702_o_0;
 wire n_8701_o_0;
 wire n_8700_o_0;
 wire n_8699_o_0;
 wire n_8698_o_0;
 wire n_8697_o_0;
 wire n_8696_o_0;
 wire n_8695_o_0;
 wire n_8694_o_0;
 wire n_8693_o_0;
 wire n_8692_o_0;
 wire n_8691_o_0;
 wire n_8690_o_0;
 wire n_8689_o_0;
 wire n_8688_o_0;
 wire n_8687_o_0;
 wire n_8686_o_0;
 wire n_8685_o_0;
 wire n_8684_o_0;
 wire n_8683_o_0;
 wire n_8682_o_0;
 wire n_8681_o_0;
 wire n_8680_o_0;
 wire n_8679_o_0;
 wire n_8678_o_0;
 wire n_8677_o_0;
 wire n_8676_o_0;
 wire n_8675_o_0;
 wire n_8674_o_0;
 wire n_8673_o_0;
 wire n_8672_o_0;
 wire n_8671_o_0;
 wire n_8670_o_0;
 wire n_8669_o_0;
 wire n_8668_o_0;
 wire n_8667_o_0;
 wire n_8666_o_0;
 wire n_8665_o_0;
 wire n_8664_o_0;
 wire n_8663_o_0;
 wire n_8662_o_0;
 wire n_8661_o_0;
 wire n_8660_o_0;
 wire n_8659_o_0;
 wire n_8658_o_0;
 wire n_8657_o_0;
 wire n_8656_o_0;
 wire n_8655_o_0;
 wire n_8654_o_0;
 wire n_8653_o_0;
 wire n_8652_o_0;
 wire n_8651_o_0;
 wire n_8650_o_0;
 wire n_8649_o_0;
 wire n_8648_o_0;
 wire n_8647_o_0;
 wire n_8646_o_0;
 wire n_8645_o_0;
 wire n_8644_o_0;
 wire n_8643_o_0;
 wire n_8642_o_0;
 wire n_8641_o_0;
 wire n_8640_o_0;
 wire n_8639_o_0;
 wire n_8638_o_0;
 wire n_8637_o_0;
 wire n_8636_o_0;
 wire n_8635_o_0;
 wire n_8634_o_0;
 wire n_8633_o_0;
 wire n_8632_o_0;
 wire n_8631_o_0;
 wire n_8630_o_0;
 wire n_8629_o_0;
 wire n_8628_o_0;
 wire n_8627_o_0;
 wire n_8626_o_0;
 wire n_8625_o_0;
 wire n_8624_o_0;
 wire n_8623_o_0;
 wire n_8622_o_0;
 wire n_8621_o_0;
 wire n_8620_o_0;
 wire n_8619_o_0;
 wire n_8618_o_0;
 wire n_8617_o_0;
 wire n_8616_o_0;
 wire n_8615_o_0;
 wire n_8614_o_0;
 wire n_8613_o_0;
 wire n_8612_o_0;
 wire n_8611_o_0;
 wire n_8610_o_0;
 wire n_8609_o_0;
 wire n_8608_o_0;
 wire n_8607_o_0;
 wire n_8606_o_0;
 wire n_8605_o_0;
 wire n_8604_o_0;
 wire n_8603_o_0;
 wire n_8602_o_0;
 wire n_8601_o_0;
 wire n_8600_o_0;
 wire n_8599_o_0;
 wire n_8598_o_0;
 wire n_8597_o_0;
 wire n_8596_o_0;
 wire n_8595_o_0;
 wire n_8594_o_0;
 wire n_8593_o_0;
 wire n_8592_o_0;
 wire n_8591_o_0;
 wire n_8590_o_0;
 wire n_8589_o_0;
 wire n_8588_o_0;
 wire n_8587_o_0;
 wire n_8586_o_0;
 wire n_8585_o_0;
 wire n_8584_o_0;
 wire n_8583_o_0;
 wire n_8582_o_0;
 wire n_8581_o_0;
 wire n_8580_o_0;
 wire n_8579_o_0;
 wire n_8578_o_0;
 wire n_8577_o_0;
 wire n_8576_o_0;
 wire n_8575_o_0;
 wire n_8574_o_0;
 wire n_8573_o_0;
 wire n_8572_o_0;
 wire n_8571_o_0;
 wire n_8570_o_0;
 wire n_8569_o_0;
 wire n_8568_o_0;
 wire n_8567_o_0;
 wire n_8566_o_0;
 wire n_8565_o_0;
 wire n_8564_o_0;
 wire n_8563_o_0;
 wire n_8562_o_0;
 wire n_8561_o_0;
 wire n_8560_o_0;
 wire n_8559_o_0;
 wire n_8558_o_0;
 wire n_8557_o_0;
 wire n_8556_o_0;
 wire n_8555_o_0;
 wire n_8554_o_0;
 wire n_8553_o_0;
 wire n_8552_o_0;
 wire n_8551_o_0;
 wire n_8550_o_0;
 wire n_8549_o_0;
 wire n_8548_o_0;
 wire n_8547_o_0;
 wire n_8546_o_0;
 wire n_8545_o_0;
 wire n_8544_o_0;
 wire n_8543_o_0;
 wire n_8542_o_0;
 wire n_8541_o_0;
 wire n_8540_o_0;
 wire n_8539_o_0;
 wire n_8538_o_0;
 wire n_8537_o_0;
 wire n_8536_o_0;
 wire n_8535_o_0;
 wire n_8534_o_0;
 wire n_8533_o_0;
 wire n_8532_o_0;
 wire n_8531_o_0;
 wire n_8530_o_0;
 wire n_8529_o_0;
 wire n_8528_o_0;
 wire n_8527_o_0;
 wire n_8526_o_0;
 wire n_8525_o_0;
 wire n_8524_o_0;
 wire n_8523_o_0;
 wire n_8522_o_0;
 wire n_8521_o_0;
 wire n_8520_o_0;
 wire n_8519_o_0;
 wire n_8518_o_0;
 wire n_8517_o_0;
 wire n_8516_o_0;
 wire n_8515_o_0;
 wire n_8514_o_0;
 wire n_8513_o_0;
 wire n_8512_o_0;
 wire n_8511_o_0;
 wire n_8510_o_0;
 wire n_8509_o_0;
 wire n_8508_o_0;
 wire n_8507_o_0;
 wire n_8506_o_0;
 wire n_8505_o_0;
 wire n_8504_o_0;
 wire n_8503_o_0;
 wire n_8502_o_0;
 wire n_8501_o_0;
 wire n_8500_o_0;
 wire n_8499_o_0;
 wire n_8498_o_0;
 wire n_8497_o_0;
 wire n_8496_o_0;
 wire n_8495_o_0;
 wire n_8494_o_0;
 wire n_8493_o_0;
 wire n_8492_o_0;
 wire n_8491_o_0;
 wire n_8490_o_0;
 wire n_8489_o_0;
 wire n_8488_o_0;
 wire n_8487_o_0;
 wire n_8486_o_0;
 wire n_8485_o_0;
 wire n_8484_o_0;
 wire n_8483_o_0;
 wire n_8482_o_0;
 wire n_8481_o_0;
 wire n_8480_o_0;
 wire n_8479_o_0;
 wire n_8478_o_0;
 wire n_8477_o_0;
 wire n_8476_o_0;
 wire n_8475_o_0;
 wire n_8474_o_0;
 wire n_8473_o_0;
 wire n_8472_o_0;
 wire n_8471_o_0;
 wire n_8470_o_0;
 wire n_8469_o_0;
 wire n_8468_o_0;
 wire n_8467_o_0;
 wire n_8466_o_0;
 wire n_8465_o_0;
 wire n_8464_o_0;
 wire n_8463_o_0;
 wire n_8462_o_0;
 wire n_8461_o_0;
 wire n_8460_o_0;
 wire n_8459_o_0;
 wire n_8458_o_0;
 wire n_8457_o_0;
 wire n_8456_o_0;
 wire n_8455_o_0;
 wire n_8454_o_0;
 wire n_8453_o_0;
 wire n_8452_o_0;
 wire n_8451_o_0;
 wire n_8450_o_0;
 wire n_8449_o_0;
 wire n_8448_o_0;
 wire n_8447_o_0;
 wire n_8446_o_0;
 wire n_8445_o_0;
 wire n_8444_o_0;
 wire n_8443_o_0;
 wire n_8442_o_0;
 wire n_8441_o_0;
 wire n_8440_o_0;
 wire n_8439_o_0;
 wire n_8438_o_0;
 wire n_8437_o_0;
 wire n_8436_o_0;
 wire n_8435_o_0;
 wire n_8434_o_0;
 wire n_8433_o_0;
 wire n_8432_o_0;
 wire n_8431_o_0;
 wire n_8430_o_0;
 wire n_8429_o_0;
 wire n_8428_o_0;
 wire n_8427_o_0;
 wire n_8426_o_0;
 wire n_8425_o_0;
 wire n_8424_o_0;
 wire n_8423_o_0;
 wire n_8422_o_0;
 wire n_8421_o_0;
 wire n_8420_o_0;
 wire n_8419_o_0;
 wire n_8418_o_0;
 wire n_8417_o_0;
 wire n_8416_o_0;
 wire n_8415_o_0;
 wire n_8414_o_0;
 wire n_8413_o_0;
 wire n_8412_o_0;
 wire n_8411_o_0;
 wire n_8410_o_0;
 wire n_8409_o_0;
 wire n_8408_o_0;
 wire n_8407_o_0;
 wire n_8406_o_0;
 wire n_8405_o_0;
 wire n_8404_o_0;
 wire n_8403_o_0;
 wire n_8402_o_0;
 wire n_8401_o_0;
 wire n_8400_o_0;
 wire n_8399_o_0;
 wire n_8398_o_0;
 wire n_8397_o_0;
 wire n_8396_o_0;
 wire n_8395_o_0;
 wire n_8394_o_0;
 wire n_8393_o_0;
 wire n_8392_o_0;
 wire n_8391_o_0;
 wire n_8390_o_0;
 wire n_8389_o_0;
 wire n_8388_o_0;
 wire n_8387_o_0;
 wire n_8386_o_0;
 wire n_8385_o_0;
 wire n_8384_o_0;
 wire n_8383_o_0;
 wire n_8382_o_0;
 wire n_8381_o_0;
 wire n_8380_o_0;
 wire n_8379_o_0;
 wire n_8378_o_0;
 wire n_8377_o_0;
 wire n_8376_o_0;
 wire n_8375_o_0;
 wire n_8374_o_0;
 wire n_8373_o_0;
 wire n_8372_o_0;
 wire n_8371_o_0;
 wire n_8370_o_0;
 wire n_8369_o_0;
 wire n_8368_o_0;
 wire n_8367_o_0;
 wire n_8366_o_0;
 wire n_8365_o_0;
 wire n_8364_o_0;
 wire n_8363_o_0;
 wire n_8362_o_0;
 wire n_8361_o_0;
 wire n_8360_o_0;
 wire n_8359_o_0;
 wire n_8358_o_0;
 wire n_8357_o_0;
 wire n_8356_o_0;
 wire n_8355_o_0;
 wire n_8354_o_0;
 wire n_8353_o_0;
 wire n_8352_o_0;
 wire n_8351_o_0;
 wire n_8350_o_0;
 wire n_8349_o_0;
 wire n_8348_o_0;
 wire n_8347_o_0;
 wire n_8346_o_0;
 wire n_8345_o_0;
 wire n_8344_o_0;
 wire n_8343_o_0;
 wire n_8342_o_0;
 wire n_8341_o_0;
 wire n_8340_o_0;
 wire n_8339_o_0;
 wire n_8338_o_0;
 wire n_8337_o_0;
 wire n_8336_o_0;
 wire n_8335_o_0;
 wire n_8334_o_0;
 wire n_8333_o_0;
 wire n_8332_o_0;
 wire n_8331_o_0;
 wire n_8330_o_0;
 wire n_8329_o_0;
 wire n_8328_o_0;
 wire n_8327_o_0;
 wire n_8326_o_0;
 wire n_8325_o_0;
 wire n_8324_o_0;
 wire n_8323_o_0;
 wire n_8322_o_0;
 wire n_8321_o_0;
 wire n_8320_o_0;
 wire n_8319_o_0;
 wire n_8318_o_0;
 wire n_8317_o_0;
 wire n_8316_o_0;
 wire n_8315_o_0;
 wire n_8314_o_0;
 wire n_8313_o_0;
 wire n_8312_o_0;
 wire n_8311_o_0;
 wire n_8310_o_0;
 wire n_8309_o_0;
 wire n_8308_o_0;
 wire n_8307_o_0;
 wire n_8306_o_0;
 wire n_8305_o_0;
 wire n_8304_o_0;
 wire n_8303_o_0;
 wire n_8302_o_0;
 wire n_8301_o_0;
 wire n_8300_o_0;
 wire n_8299_o_0;
 wire n_8298_o_0;
 wire n_8297_o_0;
 wire n_8296_o_0;
 wire n_8295_o_0;
 wire n_8294_o_0;
 wire n_8293_o_0;
 wire n_8292_o_0;
 wire n_8291_o_0;
 wire n_8290_o_0;
 wire n_8289_o_0;
 wire n_8288_o_0;
 wire n_8287_o_0;
 wire n_8286_o_0;
 wire n_8285_o_0;
 wire n_8284_o_0;
 wire n_8283_o_0;
 wire n_8282_o_0;
 wire n_8281_o_0;
 wire n_8280_o_0;
 wire n_8279_o_0;
 wire n_8278_o_0;
 wire n_8277_o_0;
 wire n_8276_o_0;
 wire n_8275_o_0;
 wire n_8274_o_0;
 wire n_8273_o_0;
 wire n_8272_o_0;
 wire n_8271_o_0;
 wire n_8270_o_0;
 wire n_8269_o_0;
 wire n_8268_o_0;
 wire n_8267_o_0;
 wire n_8266_o_0;
 wire n_8265_o_0;
 wire n_8264_o_0;
 wire n_8263_o_0;
 wire n_8262_o_0;
 wire n_8261_o_0;
 wire n_8260_o_0;
 wire n_8259_o_0;
 wire n_8258_o_0;
 wire n_8257_o_0;
 wire n_8256_o_0;
 wire n_8255_o_0;
 wire n_8254_o_0;
 wire n_8253_o_0;
 wire n_8252_o_0;
 wire n_8251_o_0;
 wire n_8250_o_0;
 wire n_8249_o_0;
 wire n_8248_o_0;
 wire n_8247_o_0;
 wire n_8246_o_0;
 wire n_8245_o_0;
 wire n_8244_o_0;
 wire n_8243_o_0;
 wire n_8242_o_0;
 wire n_8241_o_0;
 wire n_8240_o_0;
 wire n_8239_o_0;
 wire n_8238_o_0;
 wire n_8237_o_0;
 wire n_8236_o_0;
 wire n_8235_o_0;
 wire n_8234_o_0;
 wire n_8233_o_0;
 wire n_8232_o_0;
 wire n_8231_o_0;
 wire n_8230_o_0;
 wire n_8229_o_0;
 wire n_8228_o_0;
 wire n_8227_o_0;
 wire n_8226_o_0;
 wire n_8225_o_0;
 wire n_8224_o_0;
 wire n_8223_o_0;
 wire n_8222_o_0;
 wire n_8221_o_0;
 wire n_8220_o_0;
 wire n_8219_o_0;
 wire n_8218_o_0;
 wire n_8217_o_0;
 wire n_8216_o_0;
 wire n_8215_o_0;
 wire n_8214_o_0;
 wire n_8213_o_0;
 wire n_8212_o_0;
 wire n_8211_o_0;
 wire n_8210_o_0;
 wire n_8209_o_0;
 wire n_8208_o_0;
 wire n_8207_o_0;
 wire n_8206_o_0;
 wire n_8205_o_0;
 wire n_8204_o_0;
 wire n_8203_o_0;
 wire n_8202_o_0;
 wire n_8201_o_0;
 wire n_8200_o_0;
 wire n_8199_o_0;
 wire n_8198_o_0;
 wire n_8197_o_0;
 wire n_8196_o_0;
 wire n_8195_o_0;
 wire n_8194_o_0;
 wire n_8193_o_0;
 wire n_8192_o_0;
 wire n_8191_o_0;
 wire n_8190_o_0;
 wire n_8189_o_0;
 wire n_8188_o_0;
 wire n_8187_o_0;
 wire n_8186_o_0;
 wire n_8185_o_0;
 wire n_8184_o_0;
 wire n_8183_o_0;
 wire n_8182_o_0;
 wire n_8181_o_0;
 wire n_8180_o_0;
 wire n_8179_o_0;
 wire n_8178_o_0;
 wire n_8177_o_0;
 wire n_8176_o_0;
 wire n_8175_o_0;
 wire n_8174_o_0;
 wire n_8173_o_0;
 wire n_8172_o_0;
 wire n_8171_o_0;
 wire n_8170_o_0;
 wire n_8169_o_0;
 wire n_8168_o_0;
 wire n_8167_o_0;
 wire n_8166_o_0;
 wire n_8165_o_0;
 wire n_8164_o_0;
 wire n_8163_o_0;
 wire n_8162_o_0;
 wire n_8161_o_0;
 wire n_8160_o_0;
 wire n_8159_o_0;
 wire n_8158_o_0;
 wire n_8157_o_0;
 wire n_8156_o_0;
 wire n_8155_o_0;
 wire n_8154_o_0;
 wire n_8153_o_0;
 wire n_8152_o_0;
 wire n_8151_o_0;
 wire n_8150_o_0;
 wire n_8149_o_0;
 wire n_8148_o_0;
 wire n_8147_o_0;
 wire n_8146_o_0;
 wire n_8145_o_0;
 wire n_8144_o_0;
 wire n_8143_o_0;
 wire n_8142_o_0;
 wire n_8141_o_0;
 wire n_8140_o_0;
 wire n_8139_o_0;
 wire n_8138_o_0;
 wire n_8137_o_0;
 wire n_8136_o_0;
 wire n_8135_o_0;
 wire n_8134_o_0;
 wire n_8133_o_0;
 wire n_8132_o_0;
 wire n_8131_o_0;
 wire n_8130_o_0;
 wire n_8129_o_0;
 wire n_8128_o_0;
 wire n_8127_o_0;
 wire n_8126_o_0;
 wire n_8125_o_0;
 wire n_8124_o_0;
 wire n_8123_o_0;
 wire n_8122_o_0;
 wire n_8121_o_0;
 wire n_8120_o_0;
 wire n_8119_o_0;
 wire n_8118_o_0;
 wire n_8117_o_0;
 wire n_8116_o_0;
 wire n_8115_o_0;
 wire n_8114_o_0;
 wire n_8113_o_0;
 wire n_8112_o_0;
 wire n_8111_o_0;
 wire n_8110_o_0;
 wire n_8109_o_0;
 wire n_8108_o_0;
 wire n_8107_o_0;
 wire n_8106_o_0;
 wire n_8105_o_0;
 wire n_8104_o_0;
 wire n_8103_o_0;
 wire n_8102_o_0;
 wire n_8101_o_0;
 wire n_8100_o_0;
 wire n_8099_o_0;
 wire n_8098_o_0;
 wire n_8097_o_0;
 wire n_8096_o_0;
 wire n_8095_o_0;
 wire n_8094_o_0;
 wire n_8093_o_0;
 wire n_8092_o_0;
 wire n_8091_o_0;
 wire n_8090_o_0;
 wire n_8089_o_0;
 wire n_8088_o_0;
 wire n_8087_o_0;
 wire n_8086_o_0;
 wire n_8085_o_0;
 wire n_8084_o_0;
 wire n_8083_o_0;
 wire n_8082_o_0;
 wire n_8081_o_0;
 wire n_8080_o_0;
 wire n_8079_o_0;
 wire n_8078_o_0;
 wire n_8077_o_0;
 wire n_8076_o_0;
 wire n_8075_o_0;
 wire n_8074_o_0;
 wire n_8073_o_0;
 wire n_8072_o_0;
 wire n_8071_o_0;
 wire n_8070_o_0;
 wire n_8069_o_0;
 wire n_8068_o_0;
 wire n_8067_o_0;
 wire n_8066_o_0;
 wire n_8065_o_0;
 wire n_8064_o_0;
 wire n_8063_o_0;
 wire n_8062_o_0;
 wire n_8061_o_0;
 wire n_8060_o_0;
 wire n_8059_o_0;
 wire n_8058_o_0;
 wire n_8057_o_0;
 wire n_8056_o_0;
 wire n_8055_o_0;
 wire n_8054_o_0;
 wire n_8053_o_0;
 wire n_8052_o_0;
 wire n_8051_o_0;
 wire n_8050_o_0;
 wire n_8049_o_0;
 wire n_8048_o_0;
 wire n_8047_o_0;
 wire n_8046_o_0;
 wire n_8045_o_0;
 wire n_8044_o_0;
 wire n_8043_o_0;
 wire n_8042_o_0;
 wire n_8041_o_0;
 wire n_8040_o_0;
 wire n_8039_o_0;
 wire n_8038_o_0;
 wire n_8037_o_0;
 wire n_8036_o_0;
 wire n_8035_o_0;
 wire n_8034_o_0;
 wire n_8033_o_0;
 wire n_8032_o_0;
 wire n_8031_o_0;
 wire n_8030_o_0;
 wire n_8029_o_0;
 wire n_8028_o_0;
 wire n_8027_o_0;
 wire n_8026_o_0;
 wire n_8025_o_0;
 wire n_8024_o_0;
 wire n_8023_o_0;
 wire n_8022_o_0;
 wire n_8021_o_0;
 wire n_8020_o_0;
 wire n_8019_o_0;
 wire n_8018_o_0;
 wire n_8017_o_0;
 wire n_8016_o_0;
 wire n_8015_o_0;
 wire n_8014_o_0;
 wire n_8013_o_0;
 wire n_8012_o_0;
 wire n_8011_o_0;
 wire n_8010_o_0;
 wire n_8009_o_0;
 wire n_8008_o_0;
 wire n_8007_o_0;
 wire n_8006_o_0;
 wire n_8005_o_0;
 wire n_8004_o_0;
 wire n_8003_o_0;
 wire n_8002_o_0;
 wire n_8001_o_0;
 wire n_8000_o_0;
 wire n_7999_o_0;
 wire n_7998_o_0;
 wire n_7997_o_0;
 wire n_7996_o_0;
 wire n_7995_o_0;
 wire n_7994_o_0;
 wire n_7993_o_0;
 wire n_7992_o_0;
 wire n_7991_o_0;
 wire n_7990_o_0;
 wire n_7989_o_0;
 wire n_7988_o_0;
 wire n_7987_o_0;
 wire n_7986_o_0;
 wire n_7985_o_0;
 wire n_7984_o_0;
 wire n_7983_o_0;
 wire n_7982_o_0;
 wire n_7981_o_0;
 wire n_7980_o_0;
 wire n_7979_o_0;
 wire n_7978_o_0;
 wire n_7977_o_0;
 wire n_7976_o_0;
 wire n_7975_o_0;
 wire n_7974_o_0;
 wire n_7973_o_0;
 wire n_7972_o_0;
 wire n_7971_o_0;
 wire n_7970_o_0;
 wire n_7969_o_0;
 wire n_7968_o_0;
 wire n_7967_o_0;
 wire n_7966_o_0;
 wire n_7965_o_0;
 wire n_7964_o_0;
 wire n_7963_o_0;
 wire n_7962_o_0;
 wire n_7961_o_0;
 wire n_7960_o_0;
 wire n_7959_o_0;
 wire n_7958_o_0;
 wire n_7957_o_0;
 wire n_7956_o_0;
 wire n_7955_o_0;
 wire n_7954_o_0;
 wire n_7953_o_0;
 wire n_7952_o_0;
 wire n_7951_o_0;
 wire n_7950_o_0;
 wire n_7949_o_0;
 wire n_7948_o_0;
 wire n_7947_o_0;
 wire n_7946_o_0;
 wire n_7945_o_0;
 wire n_7944_o_0;
 wire n_7943_o_0;
 wire n_7942_o_0;
 wire n_7941_o_0;
 wire n_7940_o_0;
 wire n_7939_o_0;
 wire n_7938_o_0;
 wire n_7937_o_0;
 wire n_7936_o_0;
 wire n_7935_o_0;
 wire n_7934_o_0;
 wire n_7933_o_0;
 wire n_7932_o_0;
 wire n_7931_o_0;
 wire n_7930_o_0;
 wire n_7929_o_0;
 wire n_7928_o_0;
 wire n_7927_o_0;
 wire n_7926_o_0;
 wire n_7925_o_0;
 wire n_7924_o_0;
 wire n_7923_o_0;
 wire n_7922_o_0;
 wire n_7921_o_0;
 wire n_7920_o_0;
 wire n_7919_o_0;
 wire n_7918_o_0;
 wire n_7917_o_0;
 wire n_7916_o_0;
 wire n_7915_o_0;
 wire n_7914_o_0;
 wire n_7913_o_0;
 wire n_7912_o_0;
 wire n_7911_o_0;
 wire n_7910_o_0;
 wire n_7909_o_0;
 wire n_7908_o_0;
 wire n_7907_o_0;
 wire n_7906_o_0;
 wire n_7905_o_0;
 wire n_7904_o_0;
 wire n_7903_o_0;
 wire n_7902_o_0;
 wire n_7901_o_0;
 wire n_7900_o_0;
 wire n_7899_o_0;
 wire n_7898_o_0;
 wire n_7897_o_0;
 wire n_7896_o_0;
 wire n_7895_o_0;
 wire n_7894_o_0;
 wire n_7893_o_0;
 wire n_7892_o_0;
 wire n_7891_o_0;
 wire n_7890_o_0;
 wire n_7889_o_0;
 wire n_7888_o_0;
 wire n_7887_o_0;
 wire n_7886_o_0;
 wire n_7885_o_0;
 wire n_7884_o_0;
 wire n_7883_o_0;
 wire n_7882_o_0;
 wire n_7881_o_0;
 wire n_7880_o_0;
 wire n_7879_o_0;
 wire n_7878_o_0;
 wire n_7877_o_0;
 wire n_7876_o_0;
 wire n_7875_o_0;
 wire n_7874_o_0;
 wire n_7873_o_0;
 wire n_7872_o_0;
 wire n_7871_o_0;
 wire n_7870_o_0;
 wire n_7869_o_0;
 wire n_7868_o_0;
 wire n_7867_o_0;
 wire n_7866_o_0;
 wire n_7865_o_0;
 wire n_7864_o_0;
 wire n_7863_o_0;
 wire n_7862_o_0;
 wire n_7861_o_0;
 wire n_7860_o_0;
 wire n_7859_o_0;
 wire n_7858_o_0;
 wire n_7857_o_0;
 wire n_7856_o_0;
 wire n_7855_o_0;
 wire n_7854_o_0;
 wire n_7853_o_0;
 wire n_7852_o_0;
 wire n_7851_o_0;
 wire n_7850_o_0;
 wire n_7849_o_0;
 wire n_7848_o_0;
 wire n_7847_o_0;
 wire n_7846_o_0;
 wire n_7845_o_0;
 wire n_7844_o_0;
 wire n_7843_o_0;
 wire n_7842_o_0;
 wire n_7841_o_0;
 wire n_7840_o_0;
 wire n_7839_o_0;
 wire n_7838_o_0;
 wire n_7837_o_0;
 wire n_7836_o_0;
 wire n_7835_o_0;
 wire n_7834_o_0;
 wire n_7833_o_0;
 wire n_7832_o_0;
 wire n_7831_o_0;
 wire n_7830_o_0;
 wire n_7829_o_0;
 wire n_7828_o_0;
 wire n_7827_o_0;
 wire n_7826_o_0;
 wire n_7825_o_0;
 wire n_7824_o_0;
 wire n_7823_o_0;
 wire n_7822_o_0;
 wire n_7821_o_0;
 wire n_7820_o_0;
 wire n_7819_o_0;
 wire n_7818_o_0;
 wire n_7817_o_0;
 wire n_7816_o_0;
 wire n_7815_o_0;
 wire n_7814_o_0;
 wire n_7813_o_0;
 wire n_7812_o_0;
 wire n_7811_o_0;
 wire n_7810_o_0;
 wire n_7809_o_0;
 wire n_7808_o_0;
 wire n_7807_o_0;
 wire n_7806_o_0;
 wire n_7805_o_0;
 wire n_7804_o_0;
 wire n_7803_o_0;
 wire n_7802_o_0;
 wire n_7801_o_0;
 wire n_7800_o_0;
 wire n_7799_o_0;
 wire n_7798_o_0;
 wire n_7797_o_0;
 wire n_7796_o_0;
 wire n_7795_o_0;
 wire n_7794_o_0;
 wire n_7793_o_0;
 wire n_7792_o_0;
 wire n_7791_o_0;
 wire n_7790_o_0;
 wire n_7789_o_0;
 wire n_7788_o_0;
 wire n_7787_o_0;
 wire n_7786_o_0;
 wire n_7785_o_0;
 wire n_7784_o_0;
 wire n_7783_o_0;
 wire n_7782_o_0;
 wire n_7781_o_0;
 wire n_7780_o_0;
 wire n_7779_o_0;
 wire n_7778_o_0;
 wire n_7777_o_0;
 wire n_7776_o_0;
 wire n_7775_o_0;
 wire n_7774_o_0;
 wire n_7773_o_0;
 wire n_7772_o_0;
 wire n_7771_o_0;
 wire n_7770_o_0;
 wire n_7769_o_0;
 wire n_7768_o_0;
 wire n_7767_o_0;
 wire n_7766_o_0;
 wire n_7765_o_0;
 wire n_7764_o_0;
 wire n_7763_o_0;
 wire n_7762_o_0;
 wire n_7761_o_0;
 wire n_7760_o_0;
 wire n_7759_o_0;
 wire n_7758_o_0;
 wire n_7757_o_0;
 wire n_7756_o_0;
 wire n_7755_o_0;
 wire n_7754_o_0;
 wire n_7753_o_0;
 wire n_7752_o_0;
 wire n_7751_o_0;
 wire n_7750_o_0;
 wire n_7749_o_0;
 wire n_7748_o_0;
 wire n_7747_o_0;
 wire n_7746_o_0;
 wire n_7745_o_0;
 wire n_7744_o_0;
 wire n_7743_o_0;
 wire n_7742_o_0;
 wire n_7741_o_0;
 wire n_7740_o_0;
 wire n_7739_o_0;
 wire n_7738_o_0;
 wire n_7737_o_0;
 wire n_7736_o_0;
 wire n_7735_o_0;
 wire n_7734_o_0;
 wire n_7733_o_0;
 wire n_7732_o_0;
 wire n_7731_o_0;
 wire n_7730_o_0;
 wire n_7729_o_0;
 wire n_7728_o_0;
 wire n_7727_o_0;
 wire n_7726_o_0;
 wire n_7725_o_0;
 wire n_7724_o_0;
 wire n_7723_o_0;
 wire n_7722_o_0;
 wire n_7721_o_0;
 wire n_7720_o_0;
 wire n_7719_o_0;
 wire n_7718_o_0;
 wire n_7717_o_0;
 wire n_7716_o_0;
 wire n_7715_o_0;
 wire n_7714_o_0;
 wire n_7713_o_0;
 wire n_7712_o_0;
 wire n_7711_o_0;
 wire n_7710_o_0;
 wire n_7709_o_0;
 wire n_7708_o_0;
 wire n_7707_o_0;
 wire n_7706_o_0;
 wire n_7705_o_0;
 wire n_7704_o_0;
 wire n_7703_o_0;
 wire n_7702_o_0;
 wire n_7701_o_0;
 wire n_7700_o_0;
 wire n_7699_o_0;
 wire n_7698_o_0;
 wire n_7697_o_0;
 wire n_7696_o_0;
 wire n_7695_o_0;
 wire n_7694_o_0;
 wire n_7693_o_0;
 wire n_7692_o_0;
 wire n_7691_o_0;
 wire n_7690_o_0;
 wire n_7689_o_0;
 wire n_7688_o_0;
 wire n_7687_o_0;
 wire n_7686_o_0;
 wire n_7685_o_0;
 wire n_7684_o_0;
 wire n_7683_o_0;
 wire n_7682_o_0;
 wire n_7681_o_0;
 wire n_7680_o_0;
 wire n_7679_o_0;
 wire n_7678_o_0;
 wire n_7677_o_0;
 wire n_7676_o_0;
 wire n_7675_o_0;
 wire n_7674_o_0;
 wire n_7673_o_0;
 wire n_7672_o_0;
 wire n_7671_o_0;
 wire n_7670_o_0;
 wire n_7669_o_0;
 wire n_7668_o_0;
 wire n_7667_o_0;
 wire n_7666_o_0;
 wire n_7665_o_0;
 wire n_7664_o_0;
 wire n_7663_o_0;
 wire n_7662_o_0;
 wire n_7661_o_0;
 wire n_7660_o_0;
 wire n_7659_o_0;
 wire n_7658_o_0;
 wire n_7657_o_0;
 wire n_7656_o_0;
 wire n_7655_o_0;
 wire n_7654_o_0;
 wire n_7653_o_0;
 wire n_7652_o_0;
 wire n_7651_o_0;
 wire n_7650_o_0;
 wire n_7649_o_0;
 wire n_7648_o_0;
 wire n_7647_o_0;
 wire n_7646_o_0;
 wire n_7645_o_0;
 wire n_7644_o_0;
 wire n_7643_o_0;
 wire n_7642_o_0;
 wire n_7641_o_0;
 wire n_7640_o_0;
 wire n_7639_o_0;
 wire n_7638_o_0;
 wire n_7637_o_0;
 wire n_7636_o_0;
 wire n_7635_o_0;
 wire n_7634_o_0;
 wire n_7633_o_0;
 wire n_7632_o_0;
 wire n_7631_o_0;
 wire n_7630_o_0;
 wire n_7629_o_0;
 wire n_7628_o_0;
 wire n_7627_o_0;
 wire n_7626_o_0;
 wire n_7625_o_0;
 wire n_7624_o_0;
 wire n_7623_o_0;
 wire n_7622_o_0;
 wire n_7621_o_0;
 wire n_7620_o_0;
 wire n_7619_o_0;
 wire n_7618_o_0;
 wire n_7617_o_0;
 wire n_7616_o_0;
 wire n_7615_o_0;
 wire n_7614_o_0;
 wire n_7613_o_0;
 wire n_7612_o_0;
 wire n_7611_o_0;
 wire n_7610_o_0;
 wire n_7609_o_0;
 wire n_7608_o_0;
 wire n_7607_o_0;
 wire n_7606_o_0;
 wire n_7605_o_0;
 wire n_7604_o_0;
 wire n_7603_o_0;
 wire n_7602_o_0;
 wire n_7601_o_0;
 wire n_7600_o_0;
 wire n_7599_o_0;
 wire n_7598_o_0;
 wire n_7597_o_0;
 wire n_7596_o_0;
 wire n_7595_o_0;
 wire n_7594_o_0;
 wire n_7593_o_0;
 wire n_7592_o_0;
 wire n_7591_o_0;
 wire n_7590_o_0;
 wire n_7589_o_0;
 wire n_7588_o_0;
 wire n_7587_o_0;
 wire n_7586_o_0;
 wire n_7585_o_0;
 wire n_7584_o_0;
 wire n_7583_o_0;
 wire n_7582_o_0;
 wire n_7581_o_0;
 wire n_7580_o_0;
 wire n_7579_o_0;
 wire n_7578_o_0;
 wire n_7577_o_0;
 wire n_7576_o_0;
 wire n_7575_o_0;
 wire n_7574_o_0;
 wire n_7573_o_0;
 wire n_7572_o_0;
 wire n_7571_o_0;
 wire n_7570_o_0;
 wire n_7569_o_0;
 wire n_7568_o_0;
 wire n_7567_o_0;
 wire n_7566_o_0;
 wire n_7565_o_0;
 wire n_7564_o_0;
 wire n_7563_o_0;
 wire n_7562_o_0;
 wire n_7561_o_0;
 wire n_7560_o_0;
 wire n_7559_o_0;
 wire n_7558_o_0;
 wire n_7557_o_0;
 wire n_7556_o_0;
 wire n_7555_o_0;
 wire n_7554_o_0;
 wire n_7553_o_0;
 wire n_7552_o_0;
 wire n_7551_o_0;
 wire n_7550_o_0;
 wire n_7549_o_0;
 wire n_7548_o_0;
 wire n_7547_o_0;
 wire n_7546_o_0;
 wire n_7545_o_0;
 wire n_7544_o_0;
 wire n_7543_o_0;
 wire n_7542_o_0;
 wire n_7541_o_0;
 wire n_7540_o_0;
 wire n_7539_o_0;
 wire n_7538_o_0;
 wire n_7537_o_0;
 wire n_7536_o_0;
 wire n_7535_o_0;
 wire n_7534_o_0;
 wire n_7533_o_0;
 wire n_7532_o_0;
 wire n_7531_o_0;
 wire n_7530_o_0;
 wire n_7529_o_0;
 wire n_7528_o_0;
 wire n_7527_o_0;
 wire n_7526_o_0;
 wire n_7525_o_0;
 wire n_7524_o_0;
 wire n_7523_o_0;
 wire n_7522_o_0;
 wire n_7521_o_0;
 wire n_7520_o_0;
 wire n_7519_o_0;
 wire n_7518_o_0;
 wire n_7517_o_0;
 wire n_7516_o_0;
 wire n_7515_o_0;
 wire n_7514_o_0;
 wire n_7513_o_0;
 wire n_7512_o_0;
 wire n_7511_o_0;
 wire n_7510_o_0;
 wire n_7509_o_0;
 wire n_7508_o_0;
 wire n_7507_o_0;
 wire n_7506_o_0;
 wire n_7505_o_0;
 wire n_7504_o_0;
 wire n_7503_o_0;
 wire n_7502_o_0;
 wire n_7501_o_0;
 wire n_7500_o_0;
 wire n_7499_o_0;
 wire n_7498_o_0;
 wire n_7497_o_0;
 wire n_7496_o_0;
 wire n_7495_o_0;
 wire n_7494_o_0;
 wire n_7493_o_0;
 wire n_7492_o_0;
 wire n_7491_o_0;
 wire n_7490_o_0;
 wire n_7489_o_0;
 wire n_7488_o_0;
 wire n_7487_o_0;
 wire n_7486_o_0;
 wire n_7485_o_0;
 wire n_7484_o_0;
 wire n_7483_o_0;
 wire n_7482_o_0;
 wire n_7481_o_0;
 wire n_7480_o_0;
 wire n_7479_o_0;
 wire n_7478_o_0;
 wire n_7477_o_0;
 wire n_7476_o_0;
 wire n_7475_o_0;
 wire n_7474_o_0;
 wire n_7473_o_0;
 wire n_7472_o_0;
 wire n_7471_o_0;
 wire n_7470_o_0;
 wire n_7469_o_0;
 wire n_7468_o_0;
 wire n_7467_o_0;
 wire n_7466_o_0;
 wire n_7465_o_0;
 wire n_7464_o_0;
 wire n_7463_o_0;
 wire n_7462_o_0;
 wire n_7461_o_0;
 wire n_7460_o_0;
 wire n_7459_o_0;
 wire n_7458_o_0;
 wire n_7457_o_0;
 wire n_7456_o_0;
 wire n_7455_o_0;
 wire n_7454_o_0;
 wire n_7453_o_0;
 wire n_7452_o_0;
 wire n_7451_o_0;
 wire n_7450_o_0;
 wire n_7449_o_0;
 wire n_7448_o_0;
 wire n_7447_o_0;
 wire n_7446_o_0;
 wire n_7445_o_0;
 wire n_7444_o_0;
 wire n_7443_o_0;
 wire n_7442_o_0;
 wire n_7441_o_0;
 wire n_7440_o_0;
 wire n_7439_o_0;
 wire n_7438_o_0;
 wire n_7437_o_0;
 wire n_7436_o_0;
 wire n_7435_o_0;
 wire n_7434_o_0;
 wire n_7433_o_0;
 wire n_7432_o_0;
 wire n_7431_o_0;
 wire n_7430_o_0;
 wire n_7429_o_0;
 wire n_7428_o_0;
 wire n_7427_o_0;
 wire n_7426_o_0;
 wire n_7425_o_0;
 wire n_7424_o_0;
 wire n_7423_o_0;
 wire n_7422_o_0;
 wire n_7421_o_0;
 wire n_7420_o_0;
 wire n_7419_o_0;
 wire n_7418_o_0;
 wire n_7417_o_0;
 wire n_7416_o_0;
 wire n_7415_o_0;
 wire n_7414_o_0;
 wire n_7413_o_0;
 wire n_7412_o_0;
 wire n_7411_o_0;
 wire n_7410_o_0;
 wire n_7409_o_0;
 wire n_7408_o_0;
 wire n_7407_o_0;
 wire n_7406_o_0;
 wire n_7405_o_0;
 wire n_7404_o_0;
 wire n_7403_o_0;
 wire n_7402_o_0;
 wire n_7401_o_0;
 wire n_7400_o_0;
 wire n_7399_o_0;
 wire n_7398_o_0;
 wire n_7397_o_0;
 wire n_7396_o_0;
 wire n_7395_o_0;
 wire n_7394_o_0;
 wire n_7393_o_0;
 wire n_7392_o_0;
 wire n_7391_o_0;
 wire n_7390_o_0;
 wire n_7389_o_0;
 wire n_7388_o_0;
 wire n_7387_o_0;
 wire n_7386_o_0;
 wire n_7385_o_0;
 wire n_7384_o_0;
 wire n_7383_o_0;
 wire n_7382_o_0;
 wire n_7381_o_0;
 wire n_7380_o_0;
 wire n_7379_o_0;
 wire n_7378_o_0;
 wire n_7377_o_0;
 wire n_7376_o_0;
 wire n_7375_o_0;
 wire n_7374_o_0;
 wire n_7373_o_0;
 wire n_7372_o_0;
 wire n_7371_o_0;
 wire n_7370_o_0;
 wire n_7369_o_0;
 wire n_7368_o_0;
 wire n_7367_o_0;
 wire n_7366_o_0;
 wire n_7365_o_0;
 wire n_7364_o_0;
 wire n_7363_o_0;
 wire n_7362_o_0;
 wire n_7361_o_0;
 wire n_7360_o_0;
 wire n_7359_o_0;
 wire n_7358_o_0;
 wire n_7357_o_0;
 wire n_7356_o_0;
 wire n_7355_o_0;
 wire n_7354_o_0;
 wire n_7353_o_0;
 wire n_7352_o_0;
 wire n_7351_o_0;
 wire n_7350_o_0;
 wire n_7349_o_0;
 wire n_7348_o_0;
 wire n_7347_o_0;
 wire n_7346_o_0;
 wire n_7345_o_0;
 wire n_7344_o_0;
 wire n_7343_o_0;
 wire n_7342_o_0;
 wire n_7341_o_0;
 wire n_7340_o_0;
 wire n_7339_o_0;
 wire n_7338_o_0;
 wire n_7337_o_0;
 wire n_7336_o_0;
 wire n_7335_o_0;
 wire n_7334_o_0;
 wire n_7333_o_0;
 wire n_7332_o_0;
 wire n_7331_o_0;
 wire n_7330_o_0;
 wire n_7329_o_0;
 wire n_7328_o_0;
 wire n_7327_o_0;
 wire n_7326_o_0;
 wire n_7325_o_0;
 wire n_7324_o_0;
 wire n_7323_o_0;
 wire n_7322_o_0;
 wire n_7321_o_0;
 wire n_7320_o_0;
 wire n_7319_o_0;
 wire n_7318_o_0;
 wire n_7317_o_0;
 wire n_7316_o_0;
 wire n_7315_o_0;
 wire n_7314_o_0;
 wire n_7313_o_0;
 wire n_7312_o_0;
 wire n_7311_o_0;
 wire n_7310_o_0;
 wire n_7309_o_0;
 wire n_7308_o_0;
 wire n_7307_o_0;
 wire n_7306_o_0;
 wire n_7305_o_0;
 wire n_7304_o_0;
 wire n_7303_o_0;
 wire n_7302_o_0;
 wire n_7301_o_0;
 wire n_7300_o_0;
 wire n_7299_o_0;
 wire n_7298_o_0;
 wire n_7297_o_0;
 wire n_7296_o_0;
 wire n_7295_o_0;
 wire n_7294_o_0;
 wire n_7293_o_0;
 wire n_7292_o_0;
 wire n_7291_o_0;
 wire n_7290_o_0;
 wire n_7289_o_0;
 wire n_7288_o_0;
 wire n_7287_o_0;
 wire n_7286_o_0;
 wire n_7285_o_0;
 wire n_7284_o_0;
 wire n_7283_o_0;
 wire n_7282_o_0;
 wire n_7281_o_0;
 wire n_7280_o_0;
 wire n_7279_o_0;
 wire n_7278_o_0;
 wire n_7277_o_0;
 wire n_7276_o_0;
 wire n_7275_o_0;
 wire n_7274_o_0;
 wire n_7273_o_0;
 wire n_7272_o_0;
 wire n_7271_o_0;
 wire n_7270_o_0;
 wire n_7269_o_0;
 wire n_7268_o_0;
 wire n_7267_o_0;
 wire n_7266_o_0;
 wire n_7265_o_0;
 wire n_7264_o_0;
 wire n_7263_o_0;
 wire n_7262_o_0;
 wire n_7261_o_0;
 wire n_7260_o_0;
 wire n_7259_o_0;
 wire n_7258_o_0;
 wire n_7257_o_0;
 wire n_7256_o_0;
 wire n_7255_o_0;
 wire n_7254_o_0;
 wire n_7253_o_0;
 wire n_7252_o_0;
 wire n_7251_o_0;
 wire n_7250_o_0;
 wire n_7249_o_0;
 wire n_7248_o_0;
 wire n_7247_o_0;
 wire n_7246_o_0;
 wire n_7245_o_0;
 wire n_7244_o_0;
 wire n_7243_o_0;
 wire n_7242_o_0;
 wire n_7241_o_0;
 wire n_7240_o_0;
 wire n_7239_o_0;
 wire n_7238_o_0;
 wire n_7237_o_0;
 wire n_7236_o_0;
 wire n_7235_o_0;
 wire n_7234_o_0;
 wire n_7233_o_0;
 wire n_7232_o_0;
 wire n_7231_o_0;
 wire n_7230_o_0;
 wire n_7229_o_0;
 wire n_7228_o_0;
 wire n_7227_o_0;
 wire n_7226_o_0;
 wire n_7225_o_0;
 wire n_7224_o_0;
 wire n_7223_o_0;
 wire n_7222_o_0;
 wire n_7221_o_0;
 wire n_7220_o_0;
 wire n_7219_o_0;
 wire n_7218_o_0;
 wire n_7217_o_0;
 wire n_7216_o_0;
 wire n_7215_o_0;
 wire n_7214_o_0;
 wire n_7213_o_0;
 wire n_7212_o_0;
 wire n_7211_o_0;
 wire n_7210_o_0;
 wire n_7209_o_0;
 wire n_7208_o_0;
 wire n_7207_o_0;
 wire n_7206_o_0;
 wire n_7205_o_0;
 wire n_7204_o_0;
 wire n_7203_o_0;
 wire n_7202_o_0;
 wire n_7201_o_0;
 wire n_7200_o_0;
 wire n_7199_o_0;
 wire n_7198_o_0;
 wire n_7197_o_0;
 wire n_7196_o_0;
 wire n_7195_o_0;
 wire n_7194_o_0;
 wire n_7193_o_0;
 wire n_7192_o_0;
 wire n_7191_o_0;
 wire n_7190_o_0;
 wire n_7189_o_0;
 wire n_7188_o_0;
 wire n_7187_o_0;
 wire n_7186_o_0;
 wire n_7185_o_0;
 wire n_7184_o_0;
 wire n_7183_o_0;
 wire n_7182_o_0;
 wire n_7181_o_0;
 wire n_7180_o_0;
 wire n_7179_o_0;
 wire n_7178_o_0;
 wire n_7177_o_0;
 wire n_7176_o_0;
 wire n_7175_o_0;
 wire n_7174_o_0;
 wire n_7173_o_0;
 wire n_7172_o_0;
 wire n_7171_o_0;
 wire n_7170_o_0;
 wire n_7169_o_0;
 wire n_7168_o_0;
 wire n_7167_o_0;
 wire n_7166_o_0;
 wire n_7165_o_0;
 wire n_7164_o_0;
 wire n_7163_o_0;
 wire n_7162_o_0;
 wire n_7161_o_0;
 wire n_7160_o_0;
 wire n_7159_o_0;
 wire n_7158_o_0;
 wire n_7157_o_0;
 wire n_7156_o_0;
 wire n_7155_o_0;
 wire n_7154_o_0;
 wire n_7153_o_0;
 wire n_7152_o_0;
 wire n_7151_o_0;
 wire n_7150_o_0;
 wire n_7149_o_0;
 wire n_7148_o_0;
 wire n_7147_o_0;
 wire n_7146_o_0;
 wire n_7145_o_0;
 wire n_7144_o_0;
 wire n_7143_o_0;
 wire n_7142_o_0;
 wire n_7141_o_0;
 wire n_7140_o_0;
 wire n_7139_o_0;
 wire n_7138_o_0;
 wire n_7137_o_0;
 wire n_7136_o_0;
 wire n_7135_o_0;
 wire n_7134_o_0;
 wire n_7133_o_0;
 wire n_7132_o_0;
 wire n_7131_o_0;
 wire n_7130_o_0;
 wire n_7129_o_0;
 wire n_7128_o_0;
 wire n_7127_o_1;
 wire n_7127_o_0;
 wire n_7126_o_0;
 wire n_7125_o_0;
 wire n_7124_o_0;
 wire n_7123_o_0;
 wire n_7122_o_0;
 wire n_7121_o_0;
 wire n_7120_o_0;
 wire n_7119_o_0;
 wire n_7118_o_0;
 wire n_7117_o_0;
 wire n_7116_o_0;
 wire n_7115_o_0;
 wire n_7114_o_0;
 wire n_7113_o_0;
 wire n_7112_o_0;
 wire n_7111_o_0;
 wire n_7110_o_0;
 wire n_7109_o_0;
 wire n_7108_o_0;
 wire n_7107_o_0;
 wire n_7106_o_0;
 wire n_7105_o_0;
 wire n_7104_o_0;
 wire n_7103_o_0;
 wire n_7102_o_0;
 wire n_7101_o_0;
 wire n_7100_o_0;
 wire n_7099_o_0;
 wire n_7098_o_0;
 wire n_7097_o_0;
 wire n_7096_o_0;
 wire n_7095_o_0;
 wire n_7094_o_0;
 wire n_7093_o_0;
 wire n_7092_o_0;
 wire n_7091_o_0;
 wire n_7090_o_0;
 wire n_7089_o_0;
 wire n_7088_o_0;
 wire n_7087_o_0;
 wire n_7086_o_0;
 wire n_7085_o_0;
 wire n_7084_o_0;
 wire n_7083_o_0;
 wire n_7082_o_0;
 wire n_7081_o_0;
 wire n_7080_o_0;
 wire n_7079_o_0;
 wire n_7078_o_0;
 wire n_7077_o_0;
 wire n_7076_o_0;
 wire n_7075_o_0;
 wire n_7074_o_0;
 wire n_7073_o_0;
 wire n_7072_o_0;
 wire n_7071_o_0;
 wire n_7070_o_0;
 wire n_7069_o_0;
 wire n_7068_o_0;
 wire n_7067_o_0;
 wire n_7066_o_0;
 wire n_7065_o_0;
 wire n_7064_o_0;
 wire n_7063_o_0;
 wire n_7062_o_0;
 wire n_7061_o_0;
 wire n_7060_o_0;
 wire n_7059_o_0;
 wire n_7058_o_0;
 wire n_7057_o_0;
 wire n_7056_o_0;
 wire n_7055_o_0;
 wire n_7054_o_0;
 wire n_7053_o_0;
 wire n_7052_o_0;
 wire n_7051_o_0;
 wire n_7050_o_0;
 wire n_7049_o_0;
 wire n_7048_o_0;
 wire n_7047_o_0;
 wire n_7046_o_0;
 wire n_7045_o_0;
 wire n_7044_o_0;
 wire n_7043_o_0;
 wire n_7042_o_0;
 wire n_7041_o_0;
 wire n_7040_o_0;
 wire n_7039_o_0;
 wire n_7038_o_0;
 wire n_7037_o_0;
 wire n_7036_o_0;
 wire n_7035_o_0;
 wire n_7034_o_0;
 wire n_7033_o_0;
 wire n_7032_o_0;
 wire n_7031_o_0;
 wire n_7030_o_0;
 wire n_7029_o_0;
 wire n_7028_o_0;
 wire n_7027_o_0;
 wire n_7026_o_0;
 wire n_7025_o_0;
 wire n_7024_o_0;
 wire n_7023_o_0;
 wire n_7022_o_0;
 wire n_7021_o_0;
 wire n_7020_o_0;
 wire n_7019_o_0;
 wire n_7018_o_0;
 wire n_7017_o_0;
 wire n_7016_o_0;
 wire n_7015_o_0;
 wire n_7014_o_0;
 wire n_7013_o_0;
 wire n_7012_o_0;
 wire n_7011_o_0;
 wire n_7010_o_0;
 wire n_7009_o_0;
 wire n_7008_o_0;
 wire n_7007_o_0;
 wire n_7006_o_0;
 wire n_7005_o_0;
 wire n_7004_o_0;
 wire n_7003_o_0;
 wire n_7002_o_0;
 wire n_7001_o_0;
 wire n_7000_o_0;
 wire n_6999_o_0;
 wire n_6998_o_0;
 wire n_6997_o_0;
 wire n_6996_o_0;
 wire n_6995_o_0;
 wire n_6994_o_0;
 wire n_6993_o_0;
 wire n_6992_o_0;
 wire n_6991_o_0;
 wire n_6990_o_0;
 wire n_6989_o_0;
 wire n_6988_o_0;
 wire n_6987_o_0;
 wire n_6986_o_0;
 wire n_6985_o_0;
 wire n_6984_o_0;
 wire n_6983_o_0;
 wire n_6982_o_0;
 wire n_6981_o_0;
 wire n_6980_o_0;
 wire n_6979_o_0;
 wire n_6978_o_0;
 wire n_6977_o_0;
 wire n_6976_o_0;
 wire n_6975_o_0;
 wire n_6974_o_0;
 wire n_6973_o_0;
 wire n_6972_o_0;
 wire n_6971_o_0;
 wire n_6970_o_0;
 wire n_6969_o_0;
 wire n_6968_o_0;
 wire n_6967_o_0;
 wire n_6966_o_0;
 wire n_6965_o_0;
 wire n_6964_o_0;
 wire n_6963_o_0;
 wire n_6962_o_0;
 wire n_6961_o_0;
 wire n_6960_o_0;
 wire n_6959_o_0;
 wire n_6958_o_0;
 wire n_6957_o_0;
 wire n_6956_o_0;
 wire n_6955_o_0;
 wire n_6954_o_0;
 wire n_6953_o_0;
 wire n_6952_o_0;
 wire n_6951_o_0;
 wire n_6950_o_0;
 wire n_6949_o_0;
 wire n_6948_o_0;
 wire n_6947_o_0;
 wire n_6946_o_0;
 wire n_6945_o_0;
 wire n_6944_o_0;
 wire n_6943_o_0;
 wire n_6942_o_0;
 wire n_6941_o_0;
 wire n_6940_o_0;
 wire n_6939_o_0;
 wire n_6938_o_0;
 wire n_6937_o_0;
 wire n_6936_o_0;
 wire n_6935_o_0;
 wire n_6934_o_0;
 wire n_6933_o_0;
 wire n_6932_o_0;
 wire n_6931_o_0;
 wire n_6930_o_0;
 wire n_6929_o_0;
 wire n_6928_o_0;
 wire n_6927_o_0;
 wire n_6926_o_0;
 wire n_6925_o_0;
 wire n_6924_o_0;
 wire n_6923_o_0;
 wire n_6922_o_0;
 wire n_6921_o_0;
 wire n_6920_o_0;
 wire n_6919_o_0;
 wire n_6918_o_0;
 wire n_6917_o_0;
 wire n_6916_o_0;
 wire n_6915_o_0;
 wire n_6914_o_0;
 wire n_6913_o_0;
 wire n_6912_o_0;
 wire n_6911_o_0;
 wire n_6910_o_0;
 wire n_6909_o_0;
 wire n_6908_o_0;
 wire n_6907_o_0;
 wire n_6906_o_0;
 wire n_6905_o_0;
 wire n_6904_o_0;
 wire n_6903_o_0;
 wire n_6902_o_0;
 wire n_6901_o_0;
 wire n_6900_o_0;
 wire n_6899_o_0;
 wire n_6898_o_0;
 wire n_6897_o_0;
 wire n_6896_o_0;
 wire n_6895_o_0;
 wire n_6894_o_0;
 wire n_6893_o_0;
 wire n_6892_o_0;
 wire n_6891_o_0;
 wire n_6890_o_0;
 wire n_6889_o_0;
 wire n_6888_o_0;
 wire n_6887_o_0;
 wire n_6886_o_0;
 wire n_6885_o_0;
 wire n_6884_o_0;
 wire n_6883_o_0;
 wire n_6882_o_0;
 wire n_6881_o_0;
 wire n_6880_o_0;
 wire n_6879_o_0;
 wire n_6878_o_0;
 wire n_6877_o_0;
 wire n_6876_o_0;
 wire n_6875_o_0;
 wire n_6874_o_0;
 wire n_6873_o_0;
 wire n_6872_o_0;
 wire n_6871_o_0;
 wire n_6870_o_0;
 wire n_6869_o_0;
 wire n_6868_o_0;
 wire n_6867_o_0;
 wire n_6866_o_0;
 wire n_6865_o_0;
 wire n_6864_o_0;
 wire n_6863_o_0;
 wire n_6862_o_0;
 wire n_6861_o_0;
 wire n_6860_o_0;
 wire n_6859_o_0;
 wire n_6858_o_0;
 wire n_6857_o_0;
 wire n_6856_o_0;
 wire n_6855_o_1;
 wire n_6855_o_0;
 wire n_6854_o_0;
 wire n_6853_o_0;
 wire n_6852_o_0;
 wire n_6851_o_0;
 wire n_6850_o_0;
 wire n_6849_o_0;
 wire n_6848_o_0;
 wire n_6847_o_0;
 wire n_6846_o_0;
 wire n_6845_o_0;
 wire n_6844_o_0;
 wire n_6843_o_0;
 wire n_6842_o_0;
 wire n_6841_o_0;
 wire n_6840_o_0;
 wire n_6839_o_0;
 wire n_6838_o_0;
 wire n_6837_o_0;
 wire n_6836_o_0;
 wire n_6835_o_0;
 wire n_6834_o_0;
 wire n_6833_o_0;
 wire n_6832_o_0;
 wire n_6831_o_0;
 wire n_6830_o_0;
 wire n_6829_o_0;
 wire n_6828_o_0;
 wire n_6827_o_0;
 wire n_6826_o_0;
 wire n_6825_o_0;
 wire n_6824_o_0;
 wire n_6823_o_0;
 wire n_6822_o_0;
 wire n_6821_o_0;
 wire n_6820_o_0;
 wire n_6819_o_0;
 wire n_6818_o_0;
 wire n_6817_o_0;
 wire n_6816_o_0;
 wire n_6815_o_0;
 wire n_6814_o_0;
 wire n_6813_o_0;
 wire n_6812_o_0;
 wire n_6811_o_0;
 wire n_6810_o_0;
 wire n_6809_o_0;
 wire n_6808_o_0;
 wire n_6807_o_0;
 wire n_6806_o_0;
 wire n_6805_o_0;
 wire n_6804_o_0;
 wire n_6803_o_0;
 wire n_6802_o_0;
 wire n_6801_o_0;
 wire n_6800_o_0;
 wire n_6799_o_0;
 wire n_6798_o_0;
 wire n_6797_o_0;
 wire n_6796_o_0;
 wire n_6795_o_0;
 wire n_6794_o_0;
 wire n_6793_o_0;
 wire n_6792_o_0;
 wire n_6791_o_0;
 wire n_6790_o_0;
 wire n_6789_o_0;
 wire n_6788_o_0;
 wire n_6787_o_0;
 wire n_6786_o_0;
 wire n_6785_o_0;
 wire n_6784_o_0;
 wire n_6783_o_0;
 wire n_6782_o_0;
 wire n_6781_o_0;
 wire n_6780_o_0;
 wire n_6779_o_0;
 wire n_6778_o_0;
 wire n_6777_o_0;
 wire n_6776_o_0;
 wire n_6775_o_0;
 wire n_6774_o_0;
 wire n_6773_o_0;
 wire n_6772_o_0;
 wire n_6771_o_0;
 wire n_6770_o_0;
 wire n_6769_o_0;
 wire n_6768_o_0;
 wire n_6767_o_0;
 wire n_6766_o_0;
 wire n_6765_o_0;
 wire n_6764_o_0;
 wire n_6763_o_0;
 wire n_6762_o_0;
 wire n_6761_o_0;
 wire n_6760_o_0;
 wire n_6759_o_0;
 wire n_6758_o_0;
 wire n_6757_o_0;
 wire n_6756_o_0;
 wire n_6755_o_0;
 wire n_6754_o_0;
 wire n_6753_o_0;
 wire n_6752_o_0;
 wire n_6751_o_0;
 wire n_6750_o_0;
 wire n_6749_o_0;
 wire n_6748_o_0;
 wire n_6747_o_0;
 wire n_6746_o_0;
 wire n_6745_o_0;
 wire n_6744_o_0;
 wire n_6743_o_0;
 wire n_6742_o_0;
 wire n_6741_o_0;
 wire n_6740_o_0;
 wire n_6739_o_0;
 wire n_6738_o_0;
 wire n_6737_o_0;
 wire n_6736_o_0;
 wire n_6735_o_0;
 wire n_6734_o_0;
 wire n_6733_o_0;
 wire n_6732_o_0;
 wire n_6731_o_0;
 wire n_6730_o_0;
 wire n_6729_o_0;
 wire n_6728_o_0;
 wire n_6727_o_0;
 wire n_6726_o_0;
 wire n_6725_o_0;
 wire n_6724_o_0;
 wire n_6723_o_0;
 wire n_6722_o_0;
 wire n_6721_o_0;
 wire n_6720_o_0;
 wire n_6719_o_0;
 wire n_6718_o_0;
 wire n_6717_o_0;
 wire n_6716_o_0;
 wire n_6715_o_0;
 wire n_6714_o_0;
 wire n_6713_o_0;
 wire n_6712_o_0;
 wire n_6711_o_0;
 wire n_6710_o_0;
 wire n_6709_o_0;
 wire n_6708_o_0;
 wire n_6707_o_0;
 wire n_6706_o_0;
 wire n_6705_o_0;
 wire n_6704_o_0;
 wire n_6703_o_0;
 wire n_6702_o_0;
 wire n_6701_o_0;
 wire n_6700_o_0;
 wire n_6699_o_0;
 wire n_6698_o_0;
 wire n_6697_o_0;
 wire n_6696_o_0;
 wire n_6695_o_0;
 wire n_6694_o_0;
 wire n_6693_o_0;
 wire n_6692_o_0;
 wire n_6691_o_0;
 wire n_6690_o_0;
 wire n_6689_o_0;
 wire n_6688_o_0;
 wire n_6687_o_0;
 wire n_6686_o_0;
 wire n_6685_o_0;
 wire n_6684_o_0;
 wire n_6683_o_0;
 wire n_6682_o_0;
 wire n_6681_o_0;
 wire n_6680_o_0;
 wire n_6679_o_0;
 wire n_6678_o_0;
 wire n_6677_o_0;
 wire n_6676_o_0;
 wire n_6675_o_0;
 wire n_6674_o_0;
 wire n_6673_o_0;
 wire n_6672_o_0;
 wire n_6671_o_0;
 wire n_6670_o_0;
 wire n_6669_o_0;
 wire n_6668_o_0;
 wire n_6667_o_0;
 wire n_6666_o_0;
 wire n_6665_o_0;
 wire n_6664_o_0;
 wire n_6663_o_0;
 wire n_6662_o_0;
 wire n_6661_o_0;
 wire n_6660_o_0;
 wire n_6659_o_0;
 wire n_6658_o_0;
 wire n_6657_o_0;
 wire n_6656_o_0;
 wire n_6655_o_0;
 wire n_6654_o_0;
 wire n_6653_o_0;
 wire n_6652_o_0;
 wire n_6651_o_0;
 wire n_6650_o_0;
 wire n_6649_o_0;
 wire n_6648_o_0;
 wire n_6647_o_0;
 wire n_6646_o_0;
 wire n_6645_o_0;
 wire n_6644_o_0;
 wire n_6643_o_0;
 wire n_6642_o_0;
 wire n_6641_o_0;
 wire n_6640_o_0;
 wire n_6639_o_0;
 wire n_6638_o_0;
 wire n_6637_o_0;
 wire n_6636_o_0;
 wire n_6635_o_0;
 wire n_6634_o_0;
 wire n_6633_o_0;
 wire n_6632_o_0;
 wire n_6631_o_0;
 wire n_6630_o_0;
 wire n_6629_o_0;
 wire n_6628_o_0;
 wire n_6627_o_0;
 wire n_6626_o_0;
 wire n_6625_o_0;
 wire n_6624_o_0;
 wire n_6623_o_0;
 wire n_6622_o_0;
 wire n_6621_o_0;
 wire n_6620_o_0;
 wire n_6619_o_0;
 wire n_6618_o_0;
 wire n_6617_o_0;
 wire n_6616_o_0;
 wire n_6615_o_0;
 wire n_6614_o_0;
 wire n_6613_o_0;
 wire n_6612_o_0;
 wire n_6611_o_0;
 wire n_6610_o_0;
 wire n_6609_o_0;
 wire n_6608_o_0;
 wire n_6607_o_0;
 wire n_6606_o_0;
 wire n_6605_o_0;
 wire n_6604_o_0;
 wire n_6603_o_0;
 wire n_6602_o_0;
 wire n_6601_o_0;
 wire n_6600_o_0;
 wire n_6599_o_0;
 wire n_6598_o_0;
 wire n_6597_o_0;
 wire n_6596_o_0;
 wire n_6595_o_0;
 wire n_6594_o_0;
 wire n_6593_o_0;
 wire n_6592_o_0;
 wire n_6591_o_0;
 wire n_6590_o_0;
 wire n_6589_o_0;
 wire n_6588_o_0;
 wire n_6587_o_0;
 wire n_6586_o_0;
 wire n_6585_o_0;
 wire n_6584_o_0;
 wire n_6583_o_0;
 wire n_6582_o_0;
 wire n_6581_o_0;
 wire n_6580_o_0;
 wire n_6579_o_0;
 wire n_6578_o_0;
 wire n_6577_o_0;
 wire n_6576_o_0;
 wire n_6575_o_0;
 wire n_6574_o_0;
 wire n_6573_o_0;
 wire n_6572_o_0;
 wire n_6571_o_0;
 wire n_6570_o_0;
 wire n_6569_o_0;
 wire n_6568_o_0;
 wire n_6567_o_0;
 wire n_6566_o_0;
 wire n_6565_o_0;
 wire n_6564_o_0;
 wire n_6563_o_0;
 wire n_6562_o_0;
 wire n_6561_o_0;
 wire n_6560_o_0;
 wire n_6559_o_0;
 wire n_6558_o_0;
 wire n_6557_o_0;
 wire n_6556_o_0;
 wire n_6555_o_0;
 wire n_6554_o_0;
 wire n_6553_o_0;
 wire n_6552_o_0;
 wire n_6551_o_0;
 wire n_6550_o_0;
 wire n_6549_o_0;
 wire n_6548_o_0;
 wire n_6547_o_0;
 wire n_6546_o_0;
 wire n_6545_o_0;
 wire n_6544_o_0;
 wire n_6543_o_0;
 wire n_6542_o_0;
 wire n_6541_o_0;
 wire n_6540_o_0;
 wire n_6539_o_0;
 wire n_6538_o_0;
 wire n_6537_o_0;
 wire n_6536_o_0;
 wire n_6535_o_0;
 wire n_6534_o_0;
 wire n_6533_o_0;
 wire n_6532_o_0;
 wire n_6531_o_0;
 wire n_6530_o_0;
 wire n_6529_o_0;
 wire n_6528_o_0;
 wire n_6527_o_0;
 wire n_6526_o_0;
 wire n_6525_o_0;
 wire n_6524_o_0;
 wire n_6523_o_0;
 wire n_6522_o_0;
 wire n_6521_o_0;
 wire n_6520_o_0;
 wire n_6519_o_0;
 wire n_6518_o_0;
 wire n_6517_o_0;
 wire n_6516_o_0;
 wire n_6515_o_0;
 wire n_6514_o_0;
 wire n_6513_o_0;
 wire n_6512_o_0;
 wire n_6511_o_0;
 wire n_6510_o_0;
 wire n_6509_o_0;
 wire n_6508_o_0;
 wire n_6507_o_0;
 wire n_6506_o_0;
 wire n_6505_o_0;
 wire n_6504_o_0;
 wire n_6503_o_0;
 wire n_6502_o_0;
 wire n_6501_o_0;
 wire n_6500_o_0;
 wire n_6499_o_0;
 wire n_6498_o_0;
 wire n_6497_o_0;
 wire n_6496_o_0;
 wire n_6495_o_0;
 wire n_6494_o_0;
 wire n_6493_o_0;
 wire n_6492_o_0;
 wire n_6491_o_0;
 wire n_6490_o_0;
 wire n_6489_o_0;
 wire n_6488_o_0;
 wire n_6487_o_0;
 wire n_6486_o_0;
 wire n_6485_o_0;
 wire n_6484_o_0;
 wire n_6483_o_0;
 wire n_6482_o_0;
 wire n_6481_o_0;
 wire n_6480_o_0;
 wire n_6479_o_0;
 wire n_6478_o_0;
 wire n_6477_o_0;
 wire n_6476_o_0;
 wire n_6475_o_0;
 wire n_6474_o_0;
 wire n_6473_o_0;
 wire n_6472_o_0;
 wire n_6471_o_0;
 wire n_6470_o_0;
 wire n_6469_o_0;
 wire n_6468_o_0;
 wire n_6467_o_0;
 wire n_6466_o_0;
 wire n_6465_o_0;
 wire n_6464_o_0;
 wire n_6463_o_0;
 wire n_6462_o_0;
 wire n_6461_o_0;
 wire n_6460_o_0;
 wire n_6459_o_0;
 wire n_6458_o_0;
 wire n_6457_o_0;
 wire n_6456_o_0;
 wire n_6455_o_0;
 wire n_6454_o_0;
 wire n_6453_o_0;
 wire n_6452_o_0;
 wire n_6451_o_0;
 wire n_6450_o_0;
 wire n_6449_o_0;
 wire n_6448_o_0;
 wire n_6447_o_0;
 wire n_6446_o_0;
 wire n_6445_o_0;
 wire n_6444_o_0;
 wire n_6443_o_0;
 wire n_6442_o_0;
 wire n_6441_o_0;
 wire n_6440_o_0;
 wire n_6439_o_0;
 wire n_6438_o_0;
 wire n_6437_o_0;
 wire n_6436_o_0;
 wire n_6435_o_0;
 wire n_6434_o_0;
 wire n_6433_o_0;
 wire n_6432_o_0;
 wire n_6431_o_0;
 wire n_6430_o_0;
 wire n_6429_o_0;
 wire n_6428_o_0;
 wire n_6427_o_0;
 wire n_6426_o_0;
 wire n_6425_o_0;
 wire n_6424_o_0;
 wire n_6423_o_0;
 wire n_6422_o_0;
 wire n_6421_o_0;
 wire n_6420_o_0;
 wire n_6419_o_0;
 wire n_6418_o_0;
 wire n_6417_o_0;
 wire n_6416_o_0;
 wire n_6415_o_0;
 wire n_6414_o_0;
 wire n_6413_o_0;
 wire n_6412_o_0;
 wire n_6411_o_0;
 wire n_6410_o_0;
 wire n_6409_o_0;
 wire n_6408_o_0;
 wire n_6407_o_0;
 wire n_6406_o_0;
 wire n_6405_o_0;
 wire n_6404_o_0;
 wire n_6403_o_0;
 wire n_6402_o_0;
 wire n_6401_o_0;
 wire n_6400_o_0;
 wire n_6399_o_0;
 wire n_6398_o_0;
 wire n_6397_o_0;
 wire n_6396_o_0;
 wire n_6395_o_0;
 wire n_6394_o_0;
 wire n_6393_o_0;
 wire n_6392_o_0;
 wire n_6391_o_0;
 wire n_6390_o_0;
 wire n_6389_o_0;
 wire n_6388_o_0;
 wire n_6387_o_0;
 wire n_6386_o_0;
 wire n_6385_o_0;
 wire n_6384_o_0;
 wire n_6383_o_0;
 wire n_6382_o_0;
 wire n_6381_o_0;
 wire n_6380_o_0;
 wire n_6379_o_0;
 wire n_6378_o_0;
 wire n_6377_o_0;
 wire n_6376_o_0;
 wire n_6375_o_0;
 wire n_6374_o_0;
 wire n_6373_o_0;
 wire n_6372_o_0;
 wire n_6371_o_0;
 wire n_6370_o_0;
 wire n_6369_o_0;
 wire n_6368_o_0;
 wire n_6367_o_0;
 wire n_6366_o_0;
 wire n_6365_o_0;
 wire n_6364_o_0;
 wire n_6363_o_0;
 wire n_6362_o_0;
 wire n_6361_o_0;
 wire n_6360_o_0;
 wire n_6359_o_0;
 wire n_6358_o_0;
 wire n_6357_o_0;
 wire n_6356_o_0;
 wire n_6355_o_0;
 wire n_6354_o_0;
 wire n_6353_o_0;
 wire n_6352_o_0;
 wire n_6351_o_0;
 wire n_6350_o_0;
 wire n_6349_o_0;
 wire n_6348_o_0;
 wire n_6347_o_0;
 wire n_6346_o_0;
 wire n_6345_o_0;
 wire n_6344_o_0;
 wire n_6343_o_0;
 wire n_6342_o_0;
 wire n_6341_o_0;
 wire n_6340_o_0;
 wire n_6339_o_0;
 wire n_6338_o_0;
 wire n_6337_o_0;
 wire n_6336_o_0;
 wire n_6335_o_0;
 wire n_6334_o_0;
 wire n_6333_o_0;
 wire n_6332_o_0;
 wire n_6331_o_0;
 wire n_6330_o_0;
 wire n_6329_o_0;
 wire n_6328_o_0;
 wire n_6327_o_0;
 wire n_6326_o_0;
 wire n_6325_o_0;
 wire n_6324_o_0;
 wire n_6323_o_0;
 wire n_6322_o_0;
 wire n_6321_o_0;
 wire n_6320_o_0;
 wire n_6319_o_0;
 wire n_6318_o_0;
 wire n_6317_o_0;
 wire n_6316_o_0;
 wire n_6315_o_0;
 wire n_6314_o_0;
 wire n_6313_o_0;
 wire n_6312_o_0;
 wire n_6311_o_0;
 wire n_6310_o_0;
 wire n_6309_o_0;
 wire n_6308_o_0;
 wire n_6307_o_0;
 wire n_6306_o_0;
 wire n_6305_o_0;
 wire n_6304_o_0;
 wire n_6303_o_0;
 wire n_6302_o_0;
 wire n_6301_o_0;
 wire n_6300_o_0;
 wire n_6299_o_0;
 wire n_6298_o_0;
 wire n_6297_o_0;
 wire n_6296_o_0;
 wire n_6295_o_0;
 wire n_6294_o_0;
 wire n_6293_o_0;
 wire n_6292_o_0;
 wire n_6291_o_0;
 wire n_6290_o_0;
 wire n_6289_o_0;
 wire n_6288_o_0;
 wire n_6287_o_0;
 wire n_6286_o_0;
 wire n_6285_o_0;
 wire n_6284_o_0;
 wire n_6283_o_0;
 wire n_6282_o_0;
 wire n_6281_o_0;
 wire n_6280_o_0;
 wire n_6279_o_0;
 wire n_6278_o_0;
 wire n_6277_o_0;
 wire n_6276_o_0;
 wire n_6275_o_0;
 wire n_6274_o_0;
 wire n_6273_o_0;
 wire n_6272_o_0;
 wire n_6271_o_0;
 wire n_6270_o_0;
 wire n_6269_o_0;
 wire n_6268_o_0;
 wire n_6267_o_0;
 wire n_6266_o_0;
 wire n_6265_o_0;
 wire n_6264_o_0;
 wire n_6263_o_0;
 wire n_6262_o_0;
 wire n_6261_o_0;
 wire n_6260_o_0;
 wire n_6259_o_0;
 wire n_6258_o_0;
 wire n_6257_o_0;
 wire n_6256_o_0;
 wire n_6255_o_0;
 wire n_6254_o_0;
 wire n_6253_o_0;
 wire n_6252_o_0;
 wire n_6251_o_0;
 wire n_6250_o_0;
 wire n_6249_o_0;
 wire n_6248_o_0;
 wire n_6247_o_0;
 wire n_6246_o_0;
 wire n_6245_o_0;
 wire n_6244_o_0;
 wire n_6243_o_0;
 wire n_6242_o_0;
 wire n_6241_o_0;
 wire n_6240_o_0;
 wire n_6239_o_0;
 wire n_6238_o_0;
 wire n_6237_o_0;
 wire n_6236_o_0;
 wire n_6235_o_0;
 wire n_6234_o_0;
 wire n_6233_o_0;
 wire n_6232_o_0;
 wire n_6231_o_0;
 wire n_6230_o_0;
 wire n_6229_o_0;
 wire n_6228_o_0;
 wire n_6227_o_0;
 wire n_6226_o_0;
 wire n_6225_o_0;
 wire n_6224_o_0;
 wire n_6223_o_0;
 wire n_6222_o_0;
 wire n_6221_o_0;
 wire n_6220_o_0;
 wire n_6219_o_0;
 wire n_6218_o_0;
 wire n_6217_o_0;
 wire n_6216_o_0;
 wire n_6215_o_0;
 wire n_6214_o_0;
 wire n_6213_o_0;
 wire n_6212_o_0;
 wire n_6211_o_0;
 wire n_6210_o_0;
 wire n_6209_o_0;
 wire n_6208_o_0;
 wire n_6207_o_0;
 wire n_6206_o_0;
 wire n_6205_o_0;
 wire n_6204_o_0;
 wire n_6203_o_0;
 wire n_6202_o_0;
 wire n_6201_o_0;
 wire n_6200_o_0;
 wire n_6199_o_0;
 wire n_6198_o_0;
 wire n_6197_o_0;
 wire n_6196_o_0;
 wire n_6195_o_0;
 wire n_6194_o_0;
 wire n_6193_o_0;
 wire n_6192_o_0;
 wire n_6191_o_0;
 wire n_6190_o_0;
 wire n_6189_o_0;
 wire n_6188_o_0;
 wire n_6187_o_0;
 wire n_6186_o_0;
 wire n_6185_o_0;
 wire n_6184_o_0;
 wire n_6183_o_0;
 wire n_6182_o_0;
 wire n_6181_o_0;
 wire n_6180_o_0;
 wire n_6179_o_0;
 wire n_6178_o_0;
 wire n_6177_o_0;
 wire n_6176_o_0;
 wire n_6175_o_0;
 wire n_6174_o_0;
 wire n_6173_o_0;
 wire n_6172_o_0;
 wire n_6171_o_0;
 wire n_6170_o_0;
 wire n_6169_o_0;
 wire n_6168_o_0;
 wire n_6167_o_0;
 wire n_6166_o_0;
 wire n_6165_o_0;
 wire n_6164_o_0;
 wire n_6163_o_0;
 wire n_6162_o_0;
 wire n_6161_o_0;
 wire n_6160_o_0;
 wire n_6159_o_0;
 wire n_6158_o_0;
 wire n_6157_o_0;
 wire n_6156_o_0;
 wire n_6155_o_0;
 wire n_6154_o_0;
 wire n_6153_o_0;
 wire n_6152_o_0;
 wire n_6151_o_0;
 wire n_6150_o_0;
 wire n_6149_o_0;
 wire n_6148_o_0;
 wire n_6147_o_0;
 wire n_6146_o_0;
 wire n_6145_o_0;
 wire n_6144_o_0;
 wire n_6143_o_0;
 wire n_6142_o_0;
 wire n_6141_o_0;
 wire n_6140_o_0;
 wire n_6139_o_0;
 wire n_6138_o_0;
 wire n_6137_o_0;
 wire n_6136_o_0;
 wire n_6135_o_0;
 wire n_6134_o_0;
 wire n_6133_o_0;
 wire n_6132_o_0;
 wire n_6131_o_0;
 wire n_6130_o_0;
 wire n_6129_o_0;
 wire n_6128_o_0;
 wire n_6127_o_0;
 wire n_6126_o_0;
 wire n_6125_o_0;
 wire n_6124_o_0;
 wire n_6123_o_0;
 wire n_6122_o_0;
 wire n_6121_o_0;
 wire n_6120_o_0;
 wire n_6119_o_0;
 wire n_6118_o_0;
 wire n_6117_o_0;
 wire n_6116_o_0;
 wire n_6115_o_0;
 wire n_6114_o_0;
 wire n_6113_o_0;
 wire n_6112_o_0;
 wire n_6111_o_0;
 wire n_6110_o_0;
 wire n_6109_o_0;
 wire n_6108_o_0;
 wire n_6107_o_0;
 wire n_6106_o_0;
 wire n_6105_o_0;
 wire n_6104_o_0;
 wire n_6103_o_0;
 wire n_6102_o_0;
 wire n_6101_o_0;
 wire n_6100_o_0;
 wire n_6099_o_0;
 wire n_6098_o_0;
 wire n_6097_o_0;
 wire n_6096_o_0;
 wire n_6095_o_0;
 wire n_6094_o_0;
 wire n_6093_o_0;
 wire n_6092_o_0;
 wire n_6091_o_0;
 wire n_6090_o_0;
 wire n_6089_o_0;
 wire n_6088_o_0;
 wire n_6087_o_0;
 wire n_6086_o_0;
 wire n_6085_o_0;
 wire n_6084_o_0;
 wire n_6083_o_0;
 wire n_6082_o_0;
 wire n_6081_o_0;
 wire n_6080_o_0;
 wire n_6079_o_0;
 wire n_6078_o_0;
 wire n_6077_o_0;
 wire n_6076_o_0;
 wire n_6075_o_0;
 wire n_6074_o_0;
 wire n_6073_o_0;
 wire n_6072_o_0;
 wire n_6071_o_0;
 wire n_6070_o_0;
 wire n_6069_o_0;
 wire n_6068_o_0;
 wire n_6067_o_0;
 wire n_6066_o_0;
 wire n_6065_o_0;
 wire n_6064_o_0;
 wire n_6063_o_0;
 wire n_6062_o_0;
 wire n_6061_o_0;
 wire n_6060_o_0;
 wire n_6059_o_0;
 wire n_6058_o_0;
 wire n_6057_o_0;
 wire n_6056_o_0;
 wire n_6055_o_0;
 wire n_6054_o_0;
 wire n_6053_o_0;
 wire n_6052_o_0;
 wire n_6051_o_0;
 wire n_6050_o_0;
 wire n_6049_o_0;
 wire n_6048_o_0;
 wire n_6047_o_0;
 wire n_6046_o_0;
 wire n_6045_o_0;
 wire n_6044_o_0;
 wire n_6043_o_0;
 wire n_6042_o_0;
 wire n_6041_o_0;
 wire n_6040_o_0;
 wire n_6039_o_0;
 wire n_6038_o_0;
 wire n_6037_o_0;
 wire n_6036_o_0;
 wire n_6035_o_0;
 wire n_6034_o_0;
 wire n_6033_o_0;
 wire n_6032_o_0;
 wire n_6031_o_0;
 wire n_6030_o_0;
 wire n_6029_o_0;
 wire n_6028_o_0;
 wire n_6027_o_0;
 wire n_6026_o_0;
 wire n_6025_o_0;
 wire n_6024_o_0;
 wire n_6023_o_0;
 wire n_6022_o_0;
 wire n_6021_o_0;
 wire n_6020_o_0;
 wire n_6019_o_0;
 wire n_6018_o_0;
 wire n_6017_o_0;
 wire n_6016_o_0;
 wire n_6015_o_0;
 wire n_6014_o_0;
 wire n_6013_o_0;
 wire n_6012_o_0;
 wire n_6011_o_0;
 wire n_6010_o_0;
 wire n_6009_o_0;
 wire n_6008_o_0;
 wire n_6007_o_0;
 wire n_6006_o_0;
 wire n_6005_o_0;
 wire n_6004_o_0;
 wire n_6003_o_0;
 wire n_6002_o_0;
 wire n_6001_o_0;
 wire n_6000_o_0;
 wire n_5999_o_0;
 wire n_5998_o_0;
 wire n_5997_o_0;
 wire n_5996_o_0;
 wire n_5995_o_0;
 wire n_5994_o_0;
 wire n_5993_o_0;
 wire n_5992_o_0;
 wire n_5991_o_0;
 wire n_5990_o_0;
 wire n_5989_o_0;
 wire n_5988_o_0;
 wire n_5987_o_0;
 wire n_5986_o_0;
 wire n_5985_o_0;
 wire n_5984_o_0;
 wire n_5983_o_0;
 wire n_5982_o_0;
 wire n_5981_o_0;
 wire n_5980_o_0;
 wire n_5979_o_0;
 wire n_5978_o_0;
 wire n_5977_o_0;
 wire n_5976_o_0;
 wire n_5975_o_0;
 wire n_5974_o_0;
 wire n_5973_o_0;
 wire n_5972_o_0;
 wire n_5971_o_0;
 wire n_5970_o_0;
 wire n_5969_o_0;
 wire n_5968_o_0;
 wire n_5967_o_0;
 wire n_5966_o_0;
 wire n_5965_o_0;
 wire n_5964_o_0;
 wire n_5963_o_0;
 wire n_5962_o_0;
 wire n_5961_o_0;
 wire n_5960_o_0;
 wire n_5959_o_0;
 wire n_5958_o_0;
 wire n_5957_o_0;
 wire n_5956_o_0;
 wire n_5955_o_0;
 wire n_5954_o_0;
 wire n_5953_o_0;
 wire n_5952_o_0;
 wire n_5951_o_0;
 wire n_5950_o_0;
 wire n_5949_o_0;
 wire n_5948_o_0;
 wire n_5947_o_0;
 wire n_5946_o_0;
 wire n_5945_o_0;
 wire n_5944_o_0;
 wire n_5943_o_0;
 wire n_5942_o_0;
 wire n_5941_o_0;
 wire n_5940_o_0;
 wire n_5939_o_0;
 wire n_5938_o_0;
 wire n_5937_o_0;
 wire n_5936_o_0;
 wire n_5935_o_0;
 wire n_5934_o_0;
 wire n_5933_o_0;
 wire n_5932_o_0;
 wire n_5931_o_0;
 wire n_5930_o_0;
 wire n_5929_o_0;
 wire n_5928_o_0;
 wire n_5927_o_0;
 wire n_5926_o_0;
 wire n_5925_o_0;
 wire n_5924_o_0;
 wire n_5923_o_0;
 wire n_5922_o_0;
 wire n_5921_o_0;
 wire n_5920_o_0;
 wire n_5919_o_0;
 wire n_5918_o_0;
 wire n_5917_o_0;
 wire n_5916_o_0;
 wire n_5915_o_0;
 wire n_5914_o_0;
 wire n_5913_o_0;
 wire n_5912_o_0;
 wire n_5911_o_0;
 wire n_5910_o_0;
 wire n_5909_o_0;
 wire n_5908_o_0;
 wire n_5907_o_0;
 wire n_5906_o_0;
 wire n_5905_o_0;
 wire n_5904_o_0;
 wire n_5903_o_0;
 wire n_5902_o_0;
 wire n_5901_o_0;
 wire n_5900_o_0;
 wire n_5899_o_0;
 wire n_5898_o_0;
 wire n_5897_o_0;
 wire n_5896_o_0;
 wire n_5895_o_0;
 wire n_5894_o_0;
 wire n_5893_o_0;
 wire n_5892_o_0;
 wire n_5891_o_0;
 wire n_5890_o_0;
 wire n_5889_o_0;
 wire n_5888_o_0;
 wire n_5887_o_0;
 wire n_5886_o_0;
 wire n_5885_o_0;
 wire n_5884_o_0;
 wire n_5883_o_0;
 wire n_5882_o_0;
 wire n_5881_o_0;
 wire n_5880_o_0;
 wire n_5879_o_0;
 wire n_5878_o_0;
 wire n_5877_o_0;
 wire n_5876_o_0;
 wire n_5875_o_0;
 wire n_5874_o_0;
 wire n_5873_o_0;
 wire n_5872_o_0;
 wire n_5871_o_0;
 wire n_5870_o_0;
 wire n_5869_o_0;
 wire n_5868_o_0;
 wire n_5867_o_0;
 wire n_5866_o_0;
 wire n_5865_o_0;
 wire n_5864_o_0;
 wire n_5863_o_0;
 wire n_5862_o_0;
 wire n_5861_o_0;
 wire n_5860_o_0;
 wire n_5859_o_0;
 wire n_5858_o_0;
 wire n_5857_o_0;
 wire n_5856_o_0;
 wire n_5855_o_0;
 wire n_5854_o_0;
 wire n_5853_o_0;
 wire n_5852_o_0;
 wire n_5851_o_0;
 wire n_5850_o_0;
 wire n_5849_o_0;
 wire n_5848_o_0;
 wire n_5847_o_0;
 wire n_5846_o_0;
 wire n_5845_o_0;
 wire n_5844_o_0;
 wire n_5843_o_0;
 wire n_5842_o_0;
 wire n_5841_o_0;
 wire n_5840_o_0;
 wire n_5839_o_0;
 wire n_5838_o_0;
 wire n_5837_o_0;
 wire n_5836_o_0;
 wire n_5835_o_0;
 wire n_5834_o_0;
 wire n_5833_o_0;
 wire n_5832_o_0;
 wire n_5831_o_0;
 wire n_5830_o_0;
 wire n_5829_o_0;
 wire n_5828_o_0;
 wire n_5827_o_0;
 wire n_5826_o_0;
 wire n_5825_o_0;
 wire n_5824_o_0;
 wire n_5823_o_0;
 wire n_5822_o_0;
 wire n_5821_o_0;
 wire n_5820_o_0;
 wire n_5819_o_0;
 wire n_5818_o_0;
 wire n_5817_o_0;
 wire n_5816_o_0;
 wire n_5815_o_0;
 wire n_5814_o_0;
 wire n_5813_o_0;
 wire n_5812_o_0;
 wire n_5811_o_0;
 wire n_5810_o_0;
 wire n_5809_o_0;
 wire n_5808_o_0;
 wire n_5807_o_0;
 wire n_5806_o_0;
 wire n_5805_o_0;
 wire n_5804_o_0;
 wire n_5803_o_0;
 wire n_5802_o_0;
 wire n_5801_o_0;
 wire n_5800_o_0;
 wire n_5799_o_0;
 wire n_5798_o_0;
 wire n_5797_o_0;
 wire n_5796_o_0;
 wire n_5795_o_0;
 wire n_5794_o_0;
 wire n_5793_o_0;
 wire n_5792_o_0;
 wire n_5791_o_0;
 wire n_5790_o_0;
 wire n_5789_o_0;
 wire n_5788_o_0;
 wire n_5787_o_0;
 wire n_5786_o_0;
 wire n_5785_o_0;
 wire n_5784_o_0;
 wire n_5783_o_0;
 wire n_5782_o_0;
 wire n_5781_o_0;
 wire n_5780_o_0;
 wire n_5779_o_0;
 wire n_5778_o_0;
 wire n_5777_o_0;
 wire n_5776_o_0;
 wire n_5775_o_0;
 wire n_5774_o_0;
 wire n_5773_o_0;
 wire n_5772_o_0;
 wire n_5771_o_0;
 wire n_5770_o_0;
 wire n_5769_o_0;
 wire n_5768_o_0;
 wire n_5767_o_0;
 wire n_5766_o_0;
 wire n_5765_o_0;
 wire n_5764_o_0;
 wire n_5763_o_0;
 wire n_5762_o_0;
 wire n_5761_o_0;
 wire n_5760_o_0;
 wire n_5759_o_0;
 wire n_5758_o_0;
 wire n_5757_o_0;
 wire n_5756_o_0;
 wire n_5755_o_0;
 wire n_5754_o_0;
 wire n_5753_o_0;
 wire n_5752_o_0;
 wire n_5751_o_0;
 wire n_5750_o_0;
 wire n_5749_o_0;
 wire n_5748_o_0;
 wire n_5747_o_0;
 wire n_5746_o_0;
 wire n_5745_o_0;
 wire n_5744_o_0;
 wire n_5743_o_0;
 wire n_5742_o_0;
 wire n_5741_o_0;
 wire n_5740_o_0;
 wire n_5739_o_0;
 wire n_5738_o_0;
 wire n_5737_o_0;
 wire n_5736_o_0;
 wire n_5735_o_0;
 wire n_5734_o_0;
 wire n_5733_o_0;
 wire n_5732_o_0;
 wire n_5731_o_0;
 wire n_5730_o_0;
 wire n_5729_o_0;
 wire n_5728_o_0;
 wire n_5727_o_0;
 wire n_5726_o_0;
 wire n_5725_o_0;
 wire n_5724_o_0;
 wire n_5723_o_0;
 wire n_5722_o_0;
 wire n_5721_o_0;
 wire n_5720_o_0;
 wire n_5719_o_0;
 wire n_5718_o_0;
 wire n_5717_o_0;
 wire n_5716_o_0;
 wire n_5715_o_0;
 wire n_5714_o_0;
 wire n_5713_o_0;
 wire n_5712_o_0;
 wire n_5711_o_0;
 wire n_5710_o_0;
 wire n_5709_o_0;
 wire n_5708_o_0;
 wire n_5707_o_0;
 wire n_5706_o_0;
 wire n_5705_o_0;
 wire n_5704_o_0;
 wire n_5703_o_0;
 wire n_5702_o_0;
 wire n_5701_o_0;
 wire n_5700_o_0;
 wire n_5699_o_0;
 wire n_5698_o_0;
 wire n_5697_o_0;
 wire n_5696_o_0;
 wire n_5695_o_0;
 wire n_5694_o_0;
 wire n_5693_o_0;
 wire n_5692_o_0;
 wire n_5691_o_0;
 wire n_5690_o_0;
 wire n_5689_o_0;
 wire n_5688_o_0;
 wire n_5687_o_0;
 wire n_5686_o_0;
 wire n_5685_o_0;
 wire n_5684_o_0;
 wire n_5683_o_0;
 wire n_5682_o_0;
 wire n_5681_o_0;
 wire n_5680_o_0;
 wire n_5679_o_0;
 wire n_5678_o_0;
 wire n_5677_o_0;
 wire n_5676_o_0;
 wire n_5675_o_0;
 wire n_5674_o_0;
 wire n_5673_o_0;
 wire n_5672_o_0;
 wire n_5671_o_0;
 wire n_5670_o_0;
 wire n_5669_o_0;
 wire n_5668_o_0;
 wire n_5667_o_0;
 wire n_5666_o_0;
 wire n_5665_o_0;
 wire n_5664_o_0;
 wire n_5663_o_0;
 wire n_5662_o_0;
 wire n_5661_o_0;
 wire n_5660_o_0;
 wire n_5659_o_0;
 wire n_5658_o_0;
 wire n_5657_o_0;
 wire n_5656_o_0;
 wire n_5655_o_0;
 wire n_5654_o_0;
 wire n_5653_o_0;
 wire n_5652_o_0;
 wire n_5651_o_0;
 wire n_5650_o_0;
 wire n_5649_o_0;
 wire n_5648_o_0;
 wire n_5647_o_0;
 wire n_5646_o_0;
 wire n_5645_o_0;
 wire n_5644_o_0;
 wire n_5643_o_0;
 wire n_5642_o_0;
 wire n_5641_o_0;
 wire n_5640_o_0;
 wire n_5639_o_0;
 wire n_5638_o_0;
 wire n_5637_o_0;
 wire n_5636_o_0;
 wire n_5635_o_0;
 wire n_5634_o_0;
 wire n_5633_o_0;
 wire n_5632_o_0;
 wire n_5631_o_0;
 wire n_5630_o_0;
 wire n_5629_o_0;
 wire n_5628_o_0;
 wire n_5627_o_0;
 wire n_5626_o_0;
 wire n_5625_o_0;
 wire n_5624_o_0;
 wire n_5623_o_0;
 wire n_5622_o_0;
 wire n_5621_o_0;
 wire n_5620_o_0;
 wire n_5619_o_0;
 wire n_5618_o_0;
 wire n_5617_o_0;
 wire n_5616_o_0;
 wire n_5615_o_0;
 wire n_5614_o_0;
 wire n_5613_o_0;
 wire n_5612_o_0;
 wire n_5611_o_0;
 wire n_5610_o_0;
 wire n_5609_o_0;
 wire n_5608_o_0;
 wire n_5607_o_0;
 wire n_5606_o_0;
 wire n_5605_o_0;
 wire n_5604_o_0;
 wire n_5603_o_0;
 wire n_5602_o_0;
 wire n_5601_o_0;
 wire n_5600_o_0;
 wire n_5599_o_0;
 wire n_5598_o_0;
 wire n_5597_o_0;
 wire n_5596_o_0;
 wire n_5595_o_0;
 wire n_5594_o_0;
 wire n_5593_o_0;
 wire n_5592_o_0;
 wire n_5591_o_0;
 wire n_5590_o_0;
 wire n_5589_o_0;
 wire n_5588_o_0;
 wire n_5587_o_0;
 wire n_5586_o_0;
 wire n_5585_o_0;
 wire n_5584_o_0;
 wire n_5583_o_0;
 wire n_5582_o_0;
 wire n_5581_o_0;
 wire n_5580_o_0;
 wire n_5579_o_0;
 wire n_5578_o_0;
 wire n_5577_o_0;
 wire n_5576_o_0;
 wire n_5575_o_0;
 wire n_5574_o_0;
 wire n_5573_o_0;
 wire n_5572_o_0;
 wire n_5571_o_0;
 wire n_5570_o_0;
 wire n_5569_o_0;
 wire n_5568_o_0;
 wire n_5567_o_0;
 wire n_5566_o_0;
 wire n_5565_o_0;
 wire n_5564_o_0;
 wire n_5563_o_0;
 wire n_5562_o_0;
 wire n_5561_o_0;
 wire n_5560_o_0;
 wire n_5559_o_0;
 wire n_5558_o_0;
 wire n_5557_o_0;
 wire n_5556_o_0;
 wire n_5555_o_0;
 wire n_5554_o_0;
 wire n_5553_o_0;
 wire n_5552_o_0;
 wire n_5551_o_0;
 wire n_5550_o_0;
 wire n_5549_o_0;
 wire n_5548_o_0;
 wire n_5547_o_0;
 wire n_5546_o_0;
 wire n_5545_o_0;
 wire n_5544_o_0;
 wire n_5543_o_0;
 wire n_5542_o_0;
 wire n_5541_o_0;
 wire n_5540_o_0;
 wire n_5539_o_0;
 wire n_5538_o_0;
 wire n_5537_o_0;
 wire n_5536_o_0;
 wire n_5535_o_0;
 wire n_5534_o_0;
 wire n_5533_o_0;
 wire n_5532_o_0;
 wire n_5531_o_0;
 wire n_5530_o_0;
 wire n_5529_o_0;
 wire n_5528_o_0;
 wire n_5527_o_0;
 wire n_5526_o_0;
 wire n_5525_o_0;
 wire n_5524_o_0;
 wire n_5523_o_0;
 wire n_5522_o_0;
 wire n_5521_o_0;
 wire n_5520_o_0;
 wire n_5519_o_0;
 wire n_5518_o_0;
 wire n_5517_o_0;
 wire n_5516_o_0;
 wire n_5515_o_0;
 wire n_5514_o_0;
 wire n_5513_o_0;
 wire n_5512_o_0;
 wire n_5511_o_0;
 wire n_5510_o_0;
 wire n_5509_o_0;
 wire n_5508_o_0;
 wire n_5507_o_0;
 wire n_5506_o_0;
 wire n_5505_o_0;
 wire n_5504_o_0;
 wire n_5503_o_0;
 wire n_5502_o_0;
 wire n_5501_o_0;
 wire n_5500_o_0;
 wire n_5499_o_0;
 wire n_5498_o_0;
 wire n_5497_o_0;
 wire n_5496_o_0;
 wire n_5495_o_0;
 wire n_5494_o_0;
 wire n_5493_o_0;
 wire n_5492_o_0;
 wire n_5491_o_0;
 wire n_5490_o_0;
 wire n_5489_o_0;
 wire n_5488_o_0;
 wire n_5487_o_0;
 wire n_5486_o_0;
 wire n_5485_o_0;
 wire n_5484_o_0;
 wire n_5483_o_0;
 wire n_5482_o_0;
 wire n_5481_o_0;
 wire n_5480_o_0;
 wire n_5479_o_0;
 wire n_5478_o_0;
 wire n_5477_o_0;
 wire n_5476_o_0;
 wire n_5475_o_0;
 wire n_5474_o_0;
 wire n_5473_o_0;
 wire n_5472_o_0;
 wire n_5471_o_0;
 wire n_5470_o_0;
 wire n_5469_o_0;
 wire n_5468_o_0;
 wire n_5467_o_0;
 wire n_5466_o_0;
 wire n_5465_o_0;
 wire n_5464_o_0;
 wire n_5463_o_0;
 wire n_5462_o_0;
 wire n_5461_o_0;
 wire n_5460_o_0;
 wire n_5459_o_0;
 wire n_5458_o_0;
 wire n_5457_o_0;
 wire n_5456_o_0;
 wire n_5455_o_0;
 wire n_5454_o_0;
 wire n_5453_o_0;
 wire n_5452_o_0;
 wire n_5451_o_0;
 wire n_5450_o_0;
 wire n_5449_o_0;
 wire n_5448_o_0;
 wire n_5447_o_0;
 wire n_5446_o_0;
 wire n_5445_o_0;
 wire n_5444_o_0;
 wire n_5443_o_0;
 wire n_5442_o_0;
 wire n_5441_o_0;
 wire n_5440_o_0;
 wire n_5439_o_0;
 wire n_5438_o_0;
 wire n_5437_o_0;
 wire n_5436_o_0;
 wire n_5435_o_0;
 wire n_5434_o_0;
 wire n_5433_o_0;
 wire n_5432_o_0;
 wire n_5431_o_0;
 wire n_5430_o_0;
 wire n_5429_o_0;
 wire n_5428_o_0;
 wire n_5427_o_0;
 wire n_5426_o_0;
 wire n_5425_o_0;
 wire n_5424_o_0;
 wire n_5423_o_0;
 wire n_5422_o_0;
 wire n_5421_o_0;
 wire n_5420_o_0;
 wire n_5419_o_0;
 wire n_5418_o_0;
 wire n_5417_o_0;
 wire n_5416_o_0;
 wire n_5415_o_0;
 wire n_5414_o_0;
 wire n_5413_o_0;
 wire n_5412_o_0;
 wire n_5411_o_0;
 wire n_5410_o_0;
 wire n_5409_o_0;
 wire n_5408_o_0;
 wire n_5407_o_0;
 wire n_5406_o_0;
 wire n_5405_o_0;
 wire n_5404_o_0;
 wire n_5403_o_0;
 wire n_5402_o_0;
 wire n_5401_o_0;
 wire n_5400_o_0;
 wire n_5399_o_0;
 wire n_5398_o_0;
 wire n_5397_o_0;
 wire n_5396_o_0;
 wire n_5395_o_0;
 wire n_5394_o_0;
 wire n_5393_o_0;
 wire n_5392_o_0;
 wire n_5391_o_0;
 wire n_5390_o_0;
 wire n_5389_o_0;
 wire n_5388_o_0;
 wire n_5387_o_0;
 wire n_5386_o_0;
 wire n_5385_o_0;
 wire n_5384_o_0;
 wire n_5383_o_0;
 wire n_5382_o_0;
 wire n_5381_o_0;
 wire n_5380_o_0;
 wire n_5379_o_0;
 wire n_5378_o_0;
 wire n_5377_o_0;
 wire n_5376_o_0;
 wire n_5375_o_0;
 wire n_5374_o_0;
 wire n_5373_o_0;
 wire n_5372_o_0;
 wire n_5371_o_0;
 wire n_5370_o_0;
 wire n_5369_o_0;
 wire n_5368_o_0;
 wire n_5367_o_0;
 wire n_5366_o_0;
 wire n_5365_o_0;
 wire n_5364_o_0;
 wire n_5363_o_0;
 wire n_5362_o_0;
 wire n_5361_o_0;
 wire n_5360_o_0;
 wire n_5359_o_0;
 wire n_5358_o_0;
 wire n_5357_o_0;
 wire n_5356_o_0;
 wire n_5355_o_0;
 wire n_5354_o_0;
 wire n_5353_o_0;
 wire n_5352_o_0;
 wire n_5351_o_0;
 wire n_5350_o_0;
 wire n_5349_o_0;
 wire n_5348_o_0;
 wire n_5347_o_0;
 wire n_5346_o_0;
 wire n_5345_o_0;
 wire n_5344_o_0;
 wire n_5343_o_0;
 wire n_5342_o_0;
 wire n_5341_o_0;
 wire n_5340_o_0;
 wire n_5339_o_0;
 wire n_5338_o_0;
 wire n_5337_o_0;
 wire n_5336_o_0;
 wire n_5335_o_0;
 wire n_5334_o_0;
 wire n_5333_o_0;
 wire n_5332_o_0;
 wire n_5331_o_0;
 wire n_5330_o_0;
 wire n_5329_o_0;
 wire n_5328_o_0;
 wire n_5327_o_0;
 wire n_5326_o_0;
 wire n_5325_o_0;
 wire n_5324_o_0;
 wire n_5323_o_0;
 wire n_5322_o_0;
 wire n_5321_o_0;
 wire n_5320_o_0;
 wire n_5319_o_0;
 wire n_5318_o_0;
 wire n_5317_o_0;
 wire n_5316_o_0;
 wire n_5315_o_0;
 wire n_5314_o_0;
 wire n_5313_o_0;
 wire n_5312_o_0;
 wire n_5311_o_0;
 wire n_5310_o_0;
 wire n_5309_o_0;
 wire n_5308_o_0;
 wire n_5307_o_0;
 wire n_5306_o_0;
 wire n_5305_o_0;
 wire n_5304_o_0;
 wire n_5303_o_0;
 wire n_5302_o_0;
 wire n_5301_o_0;
 wire n_5300_o_0;
 wire n_5299_o_0;
 wire n_5298_o_0;
 wire n_5297_o_0;
 wire n_5296_o_0;
 wire n_5295_o_0;
 wire n_5294_o_0;
 wire n_5293_o_0;
 wire n_5292_o_0;
 wire n_5291_o_0;
 wire n_5290_o_0;
 wire n_5289_o_0;
 wire n_5288_o_0;
 wire n_5287_o_0;
 wire n_5286_o_0;
 wire n_5285_o_0;
 wire n_5284_o_0;
 wire n_5283_o_0;
 wire n_5282_o_0;
 wire n_5281_o_0;
 wire n_5280_o_0;
 wire n_5279_o_0;
 wire n_5278_o_0;
 wire n_5277_o_0;
 wire n_5276_o_0;
 wire n_5275_o_0;
 wire n_5274_o_0;
 wire n_5273_o_0;
 wire n_5272_o_0;
 wire n_5271_o_0;
 wire n_5270_o_0;
 wire n_5269_o_0;
 wire n_5268_o_0;
 wire n_5267_o_0;
 wire n_5266_o_0;
 wire n_5265_o_0;
 wire n_5264_o_0;
 wire n_5263_o_0;
 wire n_5262_o_0;
 wire n_5261_o_0;
 wire n_5260_o_0;
 wire n_5259_o_0;
 wire n_5258_o_0;
 wire n_5257_o_0;
 wire n_5256_o_0;
 wire n_5255_o_0;
 wire n_5254_o_0;
 wire n_5253_o_0;
 wire n_5252_o_0;
 wire n_5251_o_0;
 wire n_5250_o_0;
 wire n_5249_o_0;
 wire n_5248_o_0;
 wire n_5247_o_0;
 wire n_5246_o_0;
 wire n_5245_o_0;
 wire n_5244_o_0;
 wire n_5243_o_0;
 wire n_5242_o_0;
 wire n_5241_o_0;
 wire n_5240_o_0;
 wire n_5239_o_0;
 wire n_5238_o_0;
 wire n_5237_o_0;
 wire n_5236_o_0;
 wire n_5235_o_0;
 wire n_5234_o_0;
 wire n_5233_o_0;
 wire n_5232_o_0;
 wire n_5231_o_0;
 wire n_5230_o_0;
 wire n_5229_o_0;
 wire n_5228_o_0;
 wire n_5227_o_0;
 wire n_5226_o_0;
 wire n_5225_o_0;
 wire n_5224_o_0;
 wire n_5223_o_0;
 wire n_5222_o_0;
 wire n_5221_o_0;
 wire n_5220_o_0;
 wire n_5219_o_0;
 wire n_5218_o_0;
 wire n_5217_o_0;
 wire n_5216_o_0;
 wire n_5215_o_0;
 wire n_5214_o_0;
 wire n_5213_o_0;
 wire n_5212_o_0;
 wire n_5211_o_0;
 wire n_5210_o_0;
 wire n_5209_o_0;
 wire n_5208_o_0;
 wire n_5207_o_0;
 wire n_5206_o_0;
 wire n_5205_o_0;
 wire n_5204_o_0;
 wire n_5203_o_0;
 wire n_5202_o_0;
 wire n_5201_o_0;
 wire n_5200_o_0;
 wire n_5199_o_0;
 wire n_5198_o_0;
 wire n_5197_o_0;
 wire n_5196_o_0;
 wire n_5195_o_0;
 wire n_5194_o_0;
 wire n_5193_o_0;
 wire n_5192_o_0;
 wire n_5191_o_0;
 wire n_5190_o_0;
 wire n_5189_o_0;
 wire n_5188_o_0;
 wire n_5187_o_0;
 wire n_5186_o_0;
 wire n_5185_o_0;
 wire n_5184_o_0;
 wire n_5183_o_0;
 wire n_5182_o_0;
 wire n_5181_o_0;
 wire n_5180_o_0;
 wire n_5179_o_0;
 wire n_5178_o_0;
 wire n_5177_o_0;
 wire n_5176_o_0;
 wire n_5175_o_0;
 wire n_5174_o_0;
 wire n_5173_o_0;
 wire n_5172_o_0;
 wire n_5171_o_0;
 wire n_5170_o_0;
 wire n_5169_o_0;
 wire n_5168_o_0;
 wire n_5167_o_0;
 wire n_5166_o_0;
 wire n_5165_o_0;
 wire n_5164_o_0;
 wire n_5163_o_0;
 wire n_5162_o_0;
 wire n_5161_o_0;
 wire n_5160_o_0;
 wire n_5159_o_0;
 wire n_5158_o_0;
 wire n_5157_o_0;
 wire n_5156_o_0;
 wire n_5155_o_0;
 wire n_5154_o_0;
 wire n_5153_o_0;
 wire n_5152_o_0;
 wire n_5151_o_0;
 wire n_5150_o_0;
 wire n_5149_o_0;
 wire n_5148_o_0;
 wire n_5147_o_0;
 wire n_5146_o_0;
 wire n_5145_o_0;
 wire n_5144_o_0;
 wire n_5143_o_0;
 wire n_5142_o_0;
 wire n_5141_o_0;
 wire n_5140_o_0;
 wire n_5139_o_0;
 wire n_5138_o_0;
 wire n_5137_o_0;
 wire n_5136_o_0;
 wire n_5135_o_0;
 wire n_5134_o_0;
 wire n_5133_o_0;
 wire n_5132_o_0;
 wire n_5131_o_0;
 wire n_5130_o_0;
 wire n_5129_o_0;
 wire n_5128_o_0;
 wire n_5127_o_0;
 wire n_5126_o_0;
 wire n_5125_o_0;
 wire n_5124_o_0;
 wire n_5123_o_0;
 wire n_5122_o_0;
 wire n_5121_o_0;
 wire n_5120_o_0;
 wire n_5119_o_0;
 wire n_5118_o_0;
 wire n_5117_o_0;
 wire n_5116_o_0;
 wire n_5115_o_0;
 wire n_5114_o_0;
 wire n_5113_o_0;
 wire n_5112_o_0;
 wire n_5111_o_0;
 wire n_5110_o_0;
 wire n_5109_o_0;
 wire n_5108_o_0;
 wire n_5107_o_0;
 wire n_5106_o_0;
 wire n_5105_o_0;
 wire n_5104_o_0;
 wire n_5103_o_0;
 wire n_5102_o_0;
 wire n_5101_o_0;
 wire n_5100_o_0;
 wire n_5099_o_0;
 wire n_5098_o_0;
 wire n_5097_o_0;
 wire n_5096_o_0;
 wire n_5095_o_0;
 wire n_5094_o_0;
 wire n_5093_o_0;
 wire n_5092_o_0;
 wire n_5091_o_0;
 wire n_5090_o_0;
 wire n_5089_o_0;
 wire n_5088_o_0;
 wire n_5087_o_0;
 wire n_5086_o_0;
 wire n_5085_o_0;
 wire n_5084_o_0;
 wire n_5083_o_0;
 wire n_5082_o_0;
 wire n_5081_o_0;
 wire n_5080_o_0;
 wire n_5079_o_0;
 wire n_5078_o_0;
 wire n_5077_o_0;
 wire n_5076_o_0;
 wire n_5075_o_0;
 wire n_5074_o_0;
 wire n_5073_o_0;
 wire n_5072_o_0;
 wire n_5071_o_0;
 wire n_5070_o_0;
 wire n_5069_o_0;
 wire n_5068_o_0;
 wire n_5067_o_0;
 wire n_5066_o_0;
 wire n_5065_o_0;
 wire n_5064_o_0;
 wire n_5063_o_0;
 wire n_5062_o_0;
 wire n_5061_o_0;
 wire n_5060_o_0;
 wire n_5059_o_0;
 wire n_5058_o_0;
 wire n_5057_o_0;
 wire n_5056_o_0;
 wire n_5055_o_0;
 wire n_5054_o_0;
 wire n_5053_o_0;
 wire n_5052_o_0;
 wire n_5051_o_0;
 wire n_5050_o_0;
 wire n_5049_o_0;
 wire n_5048_o_0;
 wire n_5047_o_0;
 wire n_5046_o_0;
 wire n_5045_o_0;
 wire n_5044_o_0;
 wire n_5043_o_0;
 wire n_5042_o_0;
 wire n_5041_o_0;
 wire n_5040_o_0;
 wire n_5039_o_0;
 wire n_5038_o_0;
 wire n_5037_o_0;
 wire n_5036_o_0;
 wire n_5035_o_0;
 wire n_5034_o_0;
 wire n_5033_o_0;
 wire n_5032_o_0;
 wire n_5031_o_0;
 wire n_5030_o_0;
 wire n_5029_o_0;
 wire n_5028_o_0;
 wire n_5027_o_0;
 wire n_5026_o_0;
 wire n_5025_o_0;
 wire n_5024_o_0;
 wire n_5023_o_0;
 wire n_5022_o_0;
 wire n_5021_o_0;
 wire n_5020_o_0;
 wire n_5019_o_0;
 wire n_5018_o_0;
 wire n_5017_o_0;
 wire n_5016_o_0;
 wire n_5015_o_0;
 wire n_5014_o_0;
 wire n_5013_o_0;
 wire n_5012_o_0;
 wire n_5011_o_0;
 wire n_5010_o_0;
 wire n_5009_o_0;
 wire n_5008_o_0;
 wire n_5007_o_0;
 wire n_5006_o_0;
 wire n_5005_o_0;
 wire n_5004_o_0;
 wire n_5003_o_0;
 wire n_5002_o_0;
 wire n_5001_o_0;
 wire n_5000_o_0;
 wire n_4999_o_0;
 wire n_4998_o_0;
 wire n_4997_o_0;
 wire n_4996_o_0;
 wire n_4995_o_0;
 wire n_4994_o_0;
 wire n_4993_o_0;
 wire n_4992_o_0;
 wire n_4991_o_0;
 wire n_4990_o_0;
 wire n_4989_o_0;
 wire n_4988_o_0;
 wire n_4987_o_0;
 wire n_4986_o_0;
 wire n_4985_o_0;
 wire n_4984_o_0;
 wire n_4983_o_0;
 wire n_4982_o_0;
 wire n_4981_o_0;
 wire n_4980_o_0;
 wire n_4979_o_0;
 wire n_4978_o_0;
 wire n_4977_o_0;
 wire n_4976_o_0;
 wire n_4975_o_0;
 wire n_4974_o_0;
 wire n_4973_o_0;
 wire n_4972_o_0;
 wire n_4971_o_0;
 wire n_4970_o_0;
 wire n_4969_o_0;
 wire n_4968_o_0;
 wire n_4967_o_0;
 wire n_4966_o_0;
 wire n_4965_o_0;
 wire n_4964_o_0;
 wire n_4963_o_0;
 wire n_4962_o_0;
 wire n_4961_o_0;
 wire n_4960_o_0;
 wire n_4959_o_0;
 wire n_4958_o_0;
 wire n_4957_o_0;
 wire n_4956_o_0;
 wire n_4955_o_0;
 wire n_4954_o_0;
 wire n_4953_o_0;
 wire n_4952_o_0;
 wire n_4951_o_0;
 wire n_4950_o_0;
 wire n_4949_o_0;
 wire n_4948_o_0;
 wire n_4947_o_0;
 wire n_4946_o_0;
 wire n_4945_o_0;
 wire n_4944_o_0;
 wire n_4943_o_0;
 wire n_4942_o_0;
 wire n_4941_o_0;
 wire n_4940_o_0;
 wire n_4939_o_0;
 wire n_4938_o_0;
 wire n_4937_o_0;
 wire n_4936_o_0;
 wire n_4935_o_0;
 wire n_4934_o_0;
 wire n_4933_o_0;
 wire n_4932_o_0;
 wire n_4931_o_0;
 wire n_4930_o_0;
 wire n_4929_o_0;
 wire n_4928_o_0;
 wire n_4927_o_0;
 wire n_4926_o_0;
 wire n_4925_o_0;
 wire n_4924_o_0;
 wire n_4923_o_0;
 wire n_4922_o_0;
 wire n_4921_o_0;
 wire n_4920_o_0;
 wire n_4919_o_0;
 wire n_4918_o_0;
 wire n_4917_o_0;
 wire n_4916_o_0;
 wire n_4915_o_0;
 wire n_4914_o_0;
 wire n_4913_o_0;
 wire n_4912_o_0;
 wire n_4911_o_0;
 wire n_4910_o_0;
 wire n_4909_o_0;
 wire n_4908_o_0;
 wire n_4907_o_0;
 wire n_4906_o_0;
 wire n_4905_o_0;
 wire n_4904_o_0;
 wire n_4903_o_0;
 wire n_4902_o_0;
 wire n_4901_o_0;
 wire n_4900_o_0;
 wire n_4899_o_0;
 wire n_4898_o_0;
 wire n_4897_o_0;
 wire n_4896_o_0;
 wire n_4895_o_0;
 wire n_4894_o_0;
 wire n_4893_o_0;
 wire n_4892_o_0;
 wire n_4891_o_0;
 wire n_4890_o_0;
 wire n_4889_o_0;
 wire n_4888_o_0;
 wire n_4887_o_0;
 wire n_4886_o_0;
 wire n_4885_o_0;
 wire n_4884_o_0;
 wire n_4883_o_0;
 wire n_4882_o_0;
 wire n_4881_o_0;
 wire n_4880_o_0;
 wire n_4879_o_0;
 wire n_4878_o_0;
 wire n_4877_o_0;
 wire n_4876_o_0;
 wire n_4875_o_0;
 wire n_4874_o_0;
 wire n_4873_o_0;
 wire n_4872_o_0;
 wire n_4871_o_0;
 wire n_4870_o_0;
 wire n_4869_o_0;
 wire n_4868_o_0;
 wire n_4867_o_0;
 wire n_4866_o_0;
 wire n_4865_o_0;
 wire n_4864_o_0;
 wire n_4863_o_0;
 wire n_4862_o_0;
 wire n_4861_o_0;
 wire n_4860_o_0;
 wire n_4859_o_0;
 wire n_4858_o_0;
 wire n_4857_o_0;
 wire n_4856_o_0;
 wire n_4855_o_0;
 wire n_4854_o_0;
 wire n_4853_o_0;
 wire n_4852_o_0;
 wire n_4851_o_0;
 wire n_4850_o_0;
 wire n_4849_o_0;
 wire n_4848_o_0;
 wire n_4847_o_0;
 wire n_4846_o_0;
 wire n_4845_o_0;
 wire n_4844_o_0;
 wire n_4843_o_0;
 wire n_4842_o_0;
 wire n_4841_o_0;
 wire n_4840_o_0;
 wire n_4839_o_0;
 wire n_4838_o_0;
 wire n_4837_o_0;
 wire n_4836_o_0;
 wire n_4835_o_0;
 wire n_4834_o_0;
 wire n_4833_o_0;
 wire n_4832_o_0;
 wire n_4831_o_0;
 wire n_4830_o_0;
 wire n_4829_o_0;
 wire n_4828_o_0;
 wire n_4827_o_0;
 wire n_4826_o_0;
 wire n_4825_o_0;
 wire n_4824_o_0;
 wire n_4823_o_0;
 wire n_4822_o_0;
 wire n_4821_o_0;
 wire n_4820_o_0;
 wire n_4819_o_0;
 wire n_4818_o_0;
 wire n_4817_o_0;
 wire n_4816_o_0;
 wire n_4815_o_0;
 wire n_4814_o_0;
 wire n_4813_o_0;
 wire n_4812_o_0;
 wire n_4811_o_0;
 wire n_4810_o_0;
 wire n_4809_o_0;
 wire n_4808_o_0;
 wire n_4807_o_0;
 wire n_4806_o_0;
 wire n_4805_o_0;
 wire n_4804_o_0;
 wire n_4803_o_0;
 wire n_4802_o_0;
 wire n_4801_o_0;
 wire n_4800_o_0;
 wire n_4799_o_0;
 wire n_4798_o_0;
 wire n_4797_o_0;
 wire n_4796_o_0;
 wire n_4795_o_0;
 wire n_4794_o_0;
 wire n_4793_o_0;
 wire n_4792_o_0;
 wire n_4791_o_0;
 wire n_4790_o_0;
 wire n_4789_o_0;
 wire n_4788_o_0;
 wire n_4787_o_0;
 wire n_4786_o_0;
 wire n_4785_o_0;
 wire n_4784_o_0;
 wire n_4783_o_0;
 wire n_4782_o_0;
 wire n_4781_o_0;
 wire n_4780_o_0;
 wire n_4779_o_0;
 wire n_4778_o_0;
 wire n_4777_o_0;
 wire n_4776_o_0;
 wire n_4775_o_0;
 wire n_4774_o_0;
 wire n_4773_o_0;
 wire n_4772_o_0;
 wire n_4771_o_0;
 wire n_4770_o_0;
 wire n_4769_o_0;
 wire n_4768_o_0;
 wire n_4767_o_0;
 wire n_4766_o_0;
 wire n_4765_o_0;
 wire n_4764_o_0;
 wire n_4763_o_0;
 wire n_4762_o_0;
 wire n_4761_o_0;
 wire n_4760_o_0;
 wire n_4759_o_0;
 wire n_4758_o_0;
 wire n_4757_o_0;
 wire n_4756_o_0;
 wire n_4755_o_0;
 wire n_4754_o_0;
 wire n_4753_o_0;
 wire n_4752_o_0;
 wire n_4751_o_0;
 wire n_4750_o_0;
 wire n_4749_o_0;
 wire n_4748_o_0;
 wire n_4747_o_0;
 wire n_4746_o_0;
 wire n_4745_o_0;
 wire n_4744_o_0;
 wire n_4743_o_0;
 wire n_4742_o_0;
 wire n_4741_o_0;
 wire n_4740_o_0;
 wire n_4739_o_0;
 wire n_4738_o_0;
 wire n_4737_o_0;
 wire n_4736_o_0;
 wire n_4735_o_0;
 wire n_4734_o_0;
 wire n_4733_o_0;
 wire n_4732_o_0;
 wire n_4731_o_0;
 wire n_4730_o_0;
 wire n_4729_o_0;
 wire n_4728_o_0;
 wire n_4727_o_0;
 wire n_4726_o_0;
 wire n_4725_o_0;
 wire n_4724_o_0;
 wire n_4723_o_0;
 wire n_4722_o_0;
 wire n_4721_o_0;
 wire n_4720_o_0;
 wire n_4719_o_0;
 wire n_4718_o_0;
 wire n_4717_o_0;
 wire n_4716_o_0;
 wire n_4715_o_0;
 wire n_4714_o_0;
 wire n_4713_o_0;
 wire n_4712_o_0;
 wire n_4711_o_0;
 wire n_4710_o_0;
 wire n_4709_o_0;
 wire n_4708_o_0;
 wire n_4707_o_0;
 wire n_4706_o_0;
 wire n_4705_o_0;
 wire n_4704_o_0;
 wire n_4703_o_0;
 wire n_4702_o_0;
 wire n_4701_o_0;
 wire n_4700_o_0;
 wire n_4699_o_0;
 wire n_4698_o_0;
 wire n_4697_o_0;
 wire n_4696_o_0;
 wire n_4695_o_0;
 wire n_4694_o_0;
 wire n_4693_o_0;
 wire n_4692_o_0;
 wire n_4691_o_0;
 wire n_4690_o_0;
 wire n_4689_o_0;
 wire n_4688_o_0;
 wire n_4687_o_0;
 wire n_4686_o_0;
 wire n_4685_o_0;
 wire n_4684_o_0;
 wire n_4683_o_0;
 wire n_4682_o_0;
 wire n_4681_o_0;
 wire n_4680_o_0;
 wire n_4679_o_0;
 wire n_4678_o_0;
 wire n_4677_o_0;
 wire n_4676_o_0;
 wire n_4675_o_0;
 wire n_4674_o_0;
 wire n_4673_o_0;
 wire n_4672_o_0;
 wire n_4671_o_0;
 wire n_4670_o_0;
 wire n_4669_o_0;
 wire n_4668_o_0;
 wire n_4667_o_0;
 wire n_4666_o_0;
 wire n_4665_o_0;
 wire n_4664_o_0;
 wire n_4663_o_0;
 wire n_4662_o_0;
 wire n_4661_o_0;
 wire n_4660_o_0;
 wire n_4659_o_0;
 wire n_4658_o_0;
 wire n_4657_o_0;
 wire n_4656_o_0;
 wire n_4655_o_0;
 wire n_4654_o_0;
 wire n_4653_o_0;
 wire n_4652_o_0;
 wire n_4651_o_0;
 wire n_4650_o_0;
 wire n_4649_o_0;
 wire n_4648_o_0;
 wire n_4647_o_0;
 wire n_4646_o_0;
 wire n_4645_o_0;
 wire n_4644_o_0;
 wire n_4643_o_0;
 wire n_4642_o_0;
 wire n_4641_o_0;
 wire n_4640_o_0;
 wire n_4639_o_0;
 wire n_4638_o_0;
 wire n_4637_o_0;
 wire n_4636_o_0;
 wire n_4635_o_0;
 wire n_4634_o_0;
 wire n_4633_o_0;
 wire n_4632_o_0;
 wire n_4631_o_0;
 wire n_4630_o_0;
 wire n_4629_o_0;
 wire n_4628_o_0;
 wire n_4627_o_0;
 wire n_4626_o_0;
 wire n_4625_o_0;
 wire n_4624_o_0;
 wire n_4623_o_0;
 wire n_4622_o_0;
 wire n_4621_o_0;
 wire n_4620_o_0;
 wire n_4619_o_0;
 wire n_4618_o_0;
 wire n_4617_o_0;
 wire n_4616_o_0;
 wire n_4615_o_0;
 wire n_4614_o_0;
 wire n_4613_o_0;
 wire n_4612_o_0;
 wire n_4611_o_0;
 wire n_4610_o_0;
 wire n_4609_o_0;
 wire n_4608_o_0;
 wire n_4607_o_0;
 wire n_4606_o_0;
 wire n_4605_o_0;
 wire n_4604_o_0;
 wire n_4603_o_0;
 wire n_4602_o_0;
 wire n_4601_o_0;
 wire n_4600_o_0;
 wire n_4599_o_0;
 wire n_4598_o_0;
 wire n_4597_o_0;
 wire n_4596_o_0;
 wire n_4595_o_0;
 wire n_4594_o_0;
 wire n_4593_o_0;
 wire n_4592_o_0;
 wire n_4591_o_0;
 wire n_4590_o_0;
 wire n_4589_o_0;
 wire n_4588_o_0;
 wire n_4587_o_0;
 wire n_4586_o_0;
 wire n_4585_o_0;
 wire n_4584_o_0;
 wire n_4583_o_0;
 wire n_4582_o_0;
 wire n_4581_o_0;
 wire n_4580_o_0;
 wire n_4579_o_0;
 wire n_4578_o_0;
 wire n_4577_o_0;
 wire n_4576_o_0;
 wire n_4575_o_0;
 wire n_4574_o_0;
 wire n_4573_o_0;
 wire n_4572_o_0;
 wire n_4571_o_0;
 wire n_4570_o_0;
 wire n_4569_o_0;
 wire n_4568_o_0;
 wire n_4567_o_0;
 wire n_4566_o_0;
 wire n_4565_o_0;
 wire n_4564_o_0;
 wire n_4563_o_0;
 wire n_4562_o_0;
 wire n_4561_o_0;
 wire n_4560_o_0;
 wire n_4559_o_0;
 wire n_4558_o_0;
 wire n_4557_o_0;
 wire n_4556_o_0;
 wire n_4555_o_0;
 wire n_4554_o_0;
 wire n_4553_o_0;
 wire n_4552_o_0;
 wire n_4551_o_0;
 wire n_4550_o_0;
 wire n_4549_o_0;
 wire n_4548_o_0;
 wire n_4547_o_0;
 wire n_4546_o_0;
 wire n_4545_o_0;
 wire n_4544_o_0;
 wire n_4543_o_0;
 wire n_4542_o_0;
 wire n_4541_o_0;
 wire n_4540_o_0;
 wire n_4539_o_0;
 wire n_4538_o_0;
 wire n_4537_o_0;
 wire n_4536_o_0;
 wire n_4535_o_0;
 wire n_4534_o_0;
 wire n_4533_o_0;
 wire n_4532_o_0;
 wire n_4531_o_0;
 wire n_4530_o_0;
 wire n_4529_o_0;
 wire n_4528_o_0;
 wire n_4527_o_0;
 wire n_4526_o_0;
 wire n_4525_o_0;
 wire n_4524_o_0;
 wire n_4523_o_0;
 wire n_4522_o_0;
 wire n_4521_o_0;
 wire n_4520_o_0;
 wire n_4519_o_0;
 wire n_4518_o_0;
 wire n_4517_o_0;
 wire n_4516_o_0;
 wire n_4515_o_0;
 wire n_4514_o_0;
 wire n_4513_o_0;
 wire n_4512_o_0;
 wire n_4511_o_0;
 wire n_4510_o_0;
 wire n_4509_o_0;
 wire n_4508_o_0;
 wire n_4507_o_0;
 wire n_4506_o_0;
 wire n_4505_o_0;
 wire n_4504_o_0;
 wire n_4503_o_0;
 wire n_4502_o_0;
 wire n_4501_o_0;
 wire n_4500_o_0;
 wire n_4499_o_0;
 wire n_4498_o_0;
 wire n_4497_o_0;
 wire n_4496_o_0;
 wire n_4495_o_0;
 wire n_4494_o_0;
 wire n_4493_o_0;
 wire n_4492_o_0;
 wire n_4491_o_0;
 wire n_4490_o_0;
 wire n_4489_o_0;
 wire n_4488_o_0;
 wire n_4487_o_0;
 wire n_4486_o_0;
 wire n_4485_o_0;
 wire n_4484_o_0;
 wire n_4483_o_0;
 wire n_4482_o_0;
 wire n_4481_o_0;
 wire n_4480_o_0;
 wire n_4479_o_0;
 wire n_4478_o_0;
 wire n_4477_o_0;
 wire n_4476_o_0;
 wire n_4475_o_0;
 wire n_4474_o_0;
 wire n_4473_o_0;
 wire n_4472_o_0;
 wire n_4471_o_0;
 wire n_4470_o_0;
 wire n_4469_o_0;
 wire n_4468_o_0;
 wire n_4467_o_0;
 wire n_4466_o_0;
 wire n_4465_o_0;
 wire n_4464_o_0;
 wire n_4463_o_0;
 wire n_4462_o_0;
 wire n_4461_o_0;
 wire n_4460_o_0;
 wire n_4459_o_0;
 wire n_4458_o_0;
 wire n_4457_o_0;
 wire n_4456_o_0;
 wire n_4455_o_0;
 wire n_4454_o_0;
 wire n_4453_o_0;
 wire n_4452_o_0;
 wire n_4451_o_0;
 wire n_4450_o_0;
 wire n_4449_o_0;
 wire n_4448_o_0;
 wire n_4447_o_0;
 wire n_4446_o_0;
 wire n_4445_o_0;
 wire n_4444_o_0;
 wire n_4443_o_0;
 wire n_4442_o_0;
 wire n_4441_o_0;
 wire n_4440_o_0;
 wire n_4439_o_0;
 wire n_4438_o_0;
 wire n_4437_o_0;
 wire n_4436_o_0;
 wire n_4435_o_0;
 wire n_4434_o_0;
 wire n_4433_o_0;
 wire n_4432_o_0;
 wire n_4431_o_0;
 wire n_4430_o_0;
 wire n_4429_o_0;
 wire n_4428_o_0;
 wire n_4427_o_0;
 wire n_4426_o_0;
 wire n_4425_o_0;
 wire n_4424_o_0;
 wire n_4423_o_0;
 wire n_4422_o_0;
 wire n_4421_o_0;
 wire n_4420_o_0;
 wire n_4419_o_0;
 wire n_4418_o_0;
 wire n_4417_o_0;
 wire n_4416_o_0;
 wire n_4415_o_0;
 wire n_4414_o_0;
 wire n_4413_o_0;
 wire n_4412_o_0;
 wire n_4411_o_0;
 wire n_4410_o_0;
 wire n_4409_o_0;
 wire n_4408_o_0;
 wire n_4407_o_0;
 wire n_4406_o_0;
 wire n_4405_o_0;
 wire n_4404_o_0;
 wire n_4403_o_0;
 wire n_4402_o_0;
 wire n_4401_o_0;
 wire n_4400_o_0;
 wire n_4399_o_0;
 wire n_4398_o_0;
 wire n_4397_o_0;
 wire n_4396_o_0;
 wire n_4395_o_0;
 wire n_4394_o_0;
 wire n_4393_o_0;
 wire n_4392_o_0;
 wire n_4391_o_0;
 wire n_4390_o_0;
 wire n_4389_o_0;
 wire n_4388_o_0;
 wire n_4387_o_0;
 wire n_4386_o_0;
 wire n_4385_o_0;
 wire n_4384_o_0;
 wire n_4383_o_0;
 wire n_4382_o_0;
 wire n_4381_o_0;
 wire n_4380_o_0;
 wire n_4379_o_0;
 wire n_4378_o_0;
 wire n_4377_o_0;
 wire n_4376_o_0;
 wire n_4375_o_0;
 wire n_4374_o_0;
 wire n_4373_o_0;
 wire n_4372_o_0;
 wire n_4371_o_0;
 wire n_4370_o_0;
 wire n_4369_o_0;
 wire n_4368_o_0;
 wire n_4367_o_0;
 wire n_4366_o_0;
 wire n_4365_o_0;
 wire n_4364_o_0;
 wire n_4363_o_0;
 wire n_4362_o_0;
 wire n_4361_o_0;
 wire n_4360_o_0;
 wire n_4359_o_0;
 wire n_4358_o_0;
 wire n_4357_o_0;
 wire n_4356_o_0;
 wire n_4355_o_0;
 wire n_4354_o_0;
 wire n_4353_o_0;
 wire n_4352_o_0;
 wire n_4351_o_0;
 wire n_4350_o_0;
 wire n_4349_o_0;
 wire n_4348_o_0;
 wire n_4347_o_0;
 wire n_4346_o_0;
 wire n_4345_o_0;
 wire n_4344_o_0;
 wire n_4343_o_0;
 wire n_4342_o_0;
 wire n_4341_o_0;
 wire n_4340_o_0;
 wire n_4339_o_0;
 wire n_4338_o_0;
 wire n_4337_o_0;
 wire n_4336_o_0;
 wire n_4335_o_0;
 wire n_4334_o_0;
 wire n_4333_o_0;
 wire n_4332_o_0;
 wire n_4331_o_0;
 wire n_4330_o_0;
 wire n_4329_o_0;
 wire n_4328_o_0;
 wire n_4327_o_0;
 wire n_4326_o_0;
 wire n_4325_o_0;
 wire n_4324_o_0;
 wire n_4323_o_0;
 wire n_4322_o_0;
 wire n_4321_o_0;
 wire n_4320_o_0;
 wire n_4319_o_0;
 wire n_4318_o_0;
 wire n_4317_o_0;
 wire n_4316_o_0;
 wire n_4315_o_0;
 wire n_4314_o_0;
 wire n_4313_o_0;
 wire n_4312_o_0;
 wire n_4311_o_0;
 wire n_4310_o_0;
 wire n_4309_o_0;
 wire n_4308_o_0;
 wire n_4307_o_0;
 wire n_4306_o_0;
 wire n_4305_o_0;
 wire n_4304_o_0;
 wire n_4303_o_0;
 wire n_4302_o_0;
 wire n_4301_o_0;
 wire n_4300_o_0;
 wire n_4299_o_0;
 wire n_4298_o_0;
 wire n_4297_o_0;
 wire n_4296_o_0;
 wire n_4295_o_0;
 wire n_4294_o_0;
 wire n_4293_o_0;
 wire n_4292_o_0;
 wire n_4291_o_0;
 wire n_4290_o_0;
 wire n_4289_o_0;
 wire n_4288_o_0;
 wire n_4287_o_0;
 wire n_4286_o_0;
 wire n_4285_o_0;
 wire n_4284_o_0;
 wire n_4283_o_0;
 wire n_4282_o_0;
 wire n_4281_o_0;
 wire n_4280_o_0;
 wire n_4279_o_0;
 wire n_4278_o_0;
 wire n_4277_o_0;
 wire n_4276_o_0;
 wire n_4275_o_0;
 wire n_4274_o_0;
 wire n_4273_o_0;
 wire n_4272_o_0;
 wire n_4271_o_0;
 wire n_4270_o_0;
 wire n_4269_o_0;
 wire n_4268_o_0;
 wire n_4267_o_0;
 wire n_4266_o_0;
 wire n_4265_o_0;
 wire n_4264_o_0;
 wire n_4263_o_0;
 wire n_4262_o_0;
 wire n_4261_o_0;
 wire n_4260_o_0;
 wire n_4259_o_0;
 wire n_4258_o_0;
 wire n_4257_o_0;
 wire n_4256_o_0;
 wire n_4255_o_0;
 wire n_4254_o_0;
 wire n_4253_o_0;
 wire n_4252_o_0;
 wire n_4251_o_0;
 wire n_4250_o_0;
 wire n_4249_o_0;
 wire n_4248_o_0;
 wire n_4247_o_0;
 wire n_4246_o_0;
 wire n_4245_o_0;
 wire n_4244_o_0;
 wire n_4243_o_0;
 wire n_4242_o_0;
 wire n_4241_o_0;
 wire n_4240_o_0;
 wire n_4239_o_0;
 wire n_4238_o_0;
 wire n_4237_o_0;
 wire n_4236_o_0;
 wire n_4235_o_0;
 wire n_4234_o_0;
 wire n_4233_o_0;
 wire n_4232_o_0;
 wire n_4231_o_0;
 wire n_4230_o_0;
 wire n_4229_o_0;
 wire n_4228_o_0;
 wire n_4227_o_0;
 wire n_4226_o_0;
 wire n_4225_o_0;
 wire n_4224_o_0;
 wire n_4223_o_0;
 wire n_4222_o_0;
 wire n_4221_o_0;
 wire n_4220_o_0;
 wire n_4219_o_0;
 wire n_4218_o_0;
 wire n_4217_o_0;
 wire n_4216_o_0;
 wire n_4215_o_0;
 wire n_4214_o_0;
 wire n_4213_o_0;
 wire n_4212_o_0;
 wire n_4211_o_0;
 wire n_4210_o_0;
 wire n_4209_o_0;
 wire n_4208_o_0;
 wire n_4207_o_0;
 wire n_4206_o_0;
 wire n_4205_o_0;
 wire n_4204_o_0;
 wire n_4203_o_0;
 wire n_4202_o_0;
 wire n_4201_o_0;
 wire n_4200_o_0;
 wire n_4199_o_0;
 wire n_4198_o_0;
 wire n_4197_o_0;
 wire n_4196_o_0;
 wire n_4195_o_0;
 wire n_4194_o_0;
 wire n_4193_o_0;
 wire n_4192_o_0;
 wire n_4191_o_0;
 wire n_4190_o_0;
 wire n_4189_o_0;
 wire n_4188_o_0;
 wire n_4187_o_0;
 wire n_4186_o_0;
 wire n_4185_o_0;
 wire n_4184_o_0;
 wire n_4183_o_0;
 wire n_4182_o_0;
 wire n_4181_o_0;
 wire n_4180_o_0;
 wire n_4179_o_0;
 wire n_4178_o_0;
 wire n_4177_o_0;
 wire n_4176_o_0;
 wire n_4175_o_0;
 wire n_4174_o_0;
 wire n_4173_o_0;
 wire n_4172_o_0;
 wire n_4171_o_0;
 wire n_4170_o_0;
 wire n_4169_o_0;
 wire n_4168_o_0;
 wire n_4167_o_0;
 wire n_4166_o_0;
 wire n_4165_o_0;
 wire n_4164_o_0;
 wire n_4163_o_0;
 wire n_4162_o_0;
 wire n_4161_o_0;
 wire n_4160_o_0;
 wire n_4159_o_0;
 wire n_4158_o_0;
 wire n_4157_o_0;
 wire n_4156_o_0;
 wire n_4155_o_0;
 wire n_4154_o_0;
 wire n_4153_o_0;
 wire n_4152_o_0;
 wire n_4151_o_0;
 wire n_4150_o_0;
 wire n_4149_o_0;
 wire n_4148_o_0;
 wire n_4147_o_0;
 wire n_4146_o_0;
 wire n_4145_o_0;
 wire n_4144_o_0;
 wire n_4143_o_0;
 wire n_4142_o_0;
 wire n_4141_o_0;
 wire n_4140_o_0;
 wire n_4139_o_0;
 wire n_4138_o_0;
 wire n_4137_o_0;
 wire n_4136_o_0;
 wire n_4135_o_0;
 wire n_4134_o_0;
 wire n_4133_o_0;
 wire n_4132_o_0;
 wire n_4131_o_0;
 wire n_4130_o_0;
 wire n_4129_o_0;
 wire n_4128_o_0;
 wire n_4127_o_0;
 wire n_4126_o_0;
 wire n_4125_o_0;
 wire n_4124_o_0;
 wire n_4123_o_0;
 wire n_4122_o_0;
 wire n_4121_o_0;
 wire n_4120_o_0;
 wire n_4119_o_0;
 wire n_4118_o_0;
 wire n_4117_o_0;
 wire n_4116_o_0;
 wire n_4115_o_0;
 wire n_4114_o_0;
 wire n_4113_o_0;
 wire n_4112_o_0;
 wire n_4111_o_0;
 wire n_4110_o_0;
 wire n_4109_o_0;
 wire n_4108_o_0;
 wire n_4107_o_0;
 wire n_4106_o_0;
 wire n_4105_o_0;
 wire n_4104_o_0;
 wire n_4103_o_0;
 wire n_4102_o_0;
 wire n_4101_o_0;
 wire n_4100_o_0;
 wire n_4099_o_0;
 wire n_4098_o_0;
 wire n_4097_o_0;
 wire n_4096_o_0;
 wire n_4095_o_0;
 wire n_4094_o_0;
 wire n_4093_o_0;
 wire n_4092_o_0;
 wire n_4091_o_0;
 wire n_4090_o_0;
 wire n_4089_o_0;
 wire n_4088_o_0;
 wire n_4087_o_0;
 wire n_4086_o_0;
 wire n_4085_o_0;
 wire n_4084_o_0;
 wire n_4083_o_0;
 wire n_4082_o_0;
 wire n_4081_o_0;
 wire n_4080_o_0;
 wire n_4079_o_0;
 wire n_4078_o_0;
 wire n_4077_o_0;
 wire n_4076_o_0;
 wire n_4075_o_0;
 wire n_4074_o_0;
 wire n_4073_o_0;
 wire n_4072_o_0;
 wire n_4071_o_0;
 wire n_4070_o_0;
 wire n_4069_o_0;
 wire n_4068_o_0;
 wire n_4067_o_0;
 wire n_4066_o_0;
 wire n_4065_o_0;
 wire n_4064_o_0;
 wire n_4063_o_0;
 wire n_4062_o_0;
 wire n_4061_o_0;
 wire n_4060_o_0;
 wire n_4059_o_0;
 wire n_4058_o_0;
 wire n_4057_o_0;
 wire n_4056_o_0;
 wire n_4055_o_0;
 wire n_4054_o_0;
 wire n_4053_o_0;
 wire n_4052_o_0;
 wire n_4051_o_0;
 wire n_4050_o_0;
 wire n_4049_o_0;
 wire n_4048_o_0;
 wire n_4047_o_0;
 wire n_4046_o_0;
 wire n_4045_o_0;
 wire n_4044_o_0;
 wire n_4043_o_0;
 wire n_4042_o_0;
 wire n_4041_o_0;
 wire n_4040_o_0;
 wire n_4039_o_0;
 wire n_4038_o_0;
 wire n_4037_o_0;
 wire n_4036_o_0;
 wire n_4035_o_0;
 wire n_4034_o_0;
 wire n_4033_o_0;
 wire n_4032_o_0;
 wire n_4031_o_0;
 wire n_4030_o_0;
 wire n_4029_o_0;
 wire n_4028_o_0;
 wire n_4027_o_0;
 wire n_4026_o_0;
 wire n_4025_o_0;
 wire n_4024_o_0;
 wire n_4023_o_0;
 wire n_4022_o_0;
 wire n_4021_o_0;
 wire n_4020_o_0;
 wire n_4019_o_0;
 wire n_4018_o_0;
 wire n_4017_o_0;
 wire n_4016_o_0;
 wire n_4015_o_0;
 wire n_4014_o_0;
 wire n_4013_o_0;
 wire n_4012_o_0;
 wire n_4011_o_0;
 wire n_4010_o_0;
 wire n_4009_o_0;
 wire n_4008_o_0;
 wire n_4007_o_0;
 wire n_4006_o_0;
 wire n_4005_o_0;
 wire n_4004_o_0;
 wire n_4003_o_0;
 wire n_4002_o_0;
 wire n_4001_o_0;
 wire n_4000_o_0;
 wire n_3999_o_0;
 wire n_3998_o_0;
 wire n_3997_o_0;
 wire n_3996_o_0;
 wire n_3995_o_0;
 wire n_3994_o_0;
 wire n_3993_o_0;
 wire n_3992_o_0;
 wire n_3991_o_0;
 wire n_3990_o_0;
 wire n_3989_o_0;
 wire n_3988_o_0;
 wire n_3987_o_0;
 wire n_3986_o_0;
 wire n_3985_o_0;
 wire n_3984_o_0;
 wire n_3983_o_0;
 wire n_3982_o_0;
 wire n_3981_o_0;
 wire n_3980_o_0;
 wire n_3979_o_0;
 wire n_3978_o_0;
 wire n_3977_o_0;
 wire n_3976_o_0;
 wire n_3975_o_0;
 wire n_3974_o_0;
 wire n_3973_o_0;
 wire n_3972_o_0;
 wire n_3971_o_0;
 wire n_3970_o_0;
 wire n_3969_o_0;
 wire n_3968_o_0;
 wire n_3967_o_0;
 wire n_3966_o_0;
 wire n_3965_o_0;
 wire n_3964_o_0;
 wire n_3963_o_0;
 wire n_3962_o_0;
 wire n_3961_o_0;
 wire n_3960_o_0;
 wire n_3959_o_0;
 wire n_3958_o_0;
 wire n_3957_o_0;
 wire n_3956_o_0;
 wire n_3955_o_0;
 wire n_3954_o_0;
 wire n_3953_o_0;
 wire n_3952_o_0;
 wire n_3951_o_0;
 wire n_3950_o_0;
 wire n_3949_o_0;
 wire n_3948_o_0;
 wire n_3947_o_0;
 wire n_3946_o_0;
 wire n_3945_o_0;
 wire n_3944_o_0;
 wire n_3943_o_0;
 wire n_3942_o_0;
 wire n_3941_o_0;
 wire n_3940_o_0;
 wire n_3939_o_0;
 wire n_3938_o_0;
 wire n_3937_o_0;
 wire n_3936_o_0;
 wire n_3935_o_0;
 wire n_3934_o_0;
 wire n_3933_o_0;
 wire n_3932_o_0;
 wire n_3931_o_0;
 wire n_3930_o_0;
 wire n_3929_o_0;
 wire n_3928_o_0;
 wire n_3927_o_0;
 wire n_3926_o_0;
 wire n_3925_o_0;
 wire n_3924_o_0;
 wire n_3923_o_0;
 wire n_3922_o_0;
 wire n_3921_o_0;
 wire n_3920_o_0;
 wire n_3919_o_0;
 wire n_3918_o_0;
 wire n_3917_o_0;
 wire n_3916_o_0;
 wire n_3915_o_0;
 wire n_3914_o_0;
 wire n_3913_o_0;
 wire n_3912_o_0;
 wire n_3911_o_0;
 wire n_3910_o_0;
 wire n_3909_o_0;
 wire n_3908_o_0;
 wire n_3907_o_0;
 wire n_3906_o_0;
 wire n_3905_o_0;
 wire n_3904_o_0;
 wire n_3903_o_0;
 wire n_3902_o_0;
 wire n_3901_o_0;
 wire n_3900_o_0;
 wire n_3899_o_0;
 wire n_3898_o_0;
 wire n_3897_o_0;
 wire n_3896_o_0;
 wire n_3895_o_0;
 wire n_3894_o_0;
 wire n_3893_o_0;
 wire n_3892_o_0;
 wire n_3891_o_0;
 wire n_3890_o_0;
 wire n_3889_o_0;
 wire n_3888_o_0;
 wire n_3887_o_0;
 wire n_3886_o_0;
 wire n_3885_o_0;
 wire n_3884_o_0;
 wire n_3883_o_0;
 wire n_3882_o_0;
 wire n_3881_o_0;
 wire n_3880_o_0;
 wire n_3879_o_0;
 wire n_3878_o_0;
 wire n_3877_o_0;
 wire n_3876_o_0;
 wire n_3875_o_0;
 wire n_3874_o_0;
 wire n_3873_o_0;
 wire n_3872_o_0;
 wire n_3871_o_0;
 wire n_3870_o_0;
 wire n_3869_o_0;
 wire n_3868_o_0;
 wire n_3867_o_0;
 wire n_3866_o_0;
 wire n_3865_o_0;
 wire n_3864_o_0;
 wire n_3863_o_0;
 wire n_3862_o_0;
 wire n_3861_o_0;
 wire n_3860_o_0;
 wire n_3859_o_0;
 wire n_3858_o_0;
 wire n_3857_o_0;
 wire n_3856_o_0;
 wire n_3855_o_0;
 wire n_3854_o_0;
 wire n_3853_o_0;
 wire n_3852_o_0;
 wire n_3851_o_0;
 wire n_3850_o_0;
 wire n_3849_o_0;
 wire n_3848_o_0;
 wire n_3847_o_0;
 wire n_3846_o_0;
 wire n_3845_o_0;
 wire n_3844_o_0;
 wire n_3843_o_0;
 wire n_3842_o_0;
 wire n_3841_o_0;
 wire n_3840_o_0;
 wire n_3839_o_0;
 wire n_3838_o_0;
 wire n_3837_o_0;
 wire n_3836_o_0;
 wire n_3835_o_0;
 wire n_3834_o_0;
 wire n_3833_o_0;
 wire n_3832_o_0;
 wire n_3831_o_0;
 wire n_3830_o_0;
 wire n_3829_o_0;
 wire n_3828_o_0;
 wire n_3827_o_0;
 wire n_3826_o_0;
 wire n_3825_o_0;
 wire n_3824_o_0;
 wire n_3823_o_0;
 wire n_3822_o_0;
 wire n_3821_o_0;
 wire n_3820_o_0;
 wire n_3819_o_0;
 wire n_3818_o_0;
 wire n_3817_o_0;
 wire n_3816_o_0;
 wire n_3815_o_0;
 wire n_3814_o_0;
 wire n_3813_o_0;
 wire n_3812_o_0;
 wire n_3811_o_0;
 wire n_3810_o_0;
 wire n_3809_o_0;
 wire n_3808_o_0;
 wire n_3807_o_0;
 wire n_3806_o_0;
 wire n_3805_o_0;
 wire n_3804_o_0;
 wire n_3803_o_0;
 wire n_3802_o_0;
 wire n_3801_o_0;
 wire n_3800_o_0;
 wire n_3799_o_0;
 wire n_3798_o_0;
 wire n_3797_o_0;
 wire n_3796_o_0;
 wire n_3795_o_0;
 wire n_3794_o_0;
 wire n_3793_o_0;
 wire n_3792_o_0;
 wire n_3791_o_0;
 wire n_3790_o_0;
 wire n_3789_o_0;
 wire n_3788_o_0;
 wire n_3787_o_0;
 wire n_3786_o_0;
 wire n_3785_o_0;
 wire n_3784_o_0;
 wire n_3783_o_0;
 wire n_3782_o_0;
 wire n_3781_o_0;
 wire n_3780_o_0;
 wire n_3779_o_0;
 wire n_3778_o_0;
 wire n_3777_o_0;
 wire n_3776_o_0;
 wire n_3775_o_0;
 wire n_3774_o_0;
 wire n_3773_o_0;
 wire n_3772_o_0;
 wire n_3771_o_0;
 wire n_3770_o_0;
 wire n_3769_o_0;
 wire n_3768_o_0;
 wire n_3767_o_0;
 wire n_3766_o_0;
 wire n_3765_o_0;
 wire n_3764_o_0;
 wire n_3763_o_0;
 wire n_3762_o_0;
 wire n_3761_o_0;
 wire n_3760_o_0;
 wire n_3759_o_0;
 wire n_3758_o_0;
 wire n_3757_o_0;
 wire n_3756_o_0;
 wire n_3755_o_0;
 wire n_3754_o_0;
 wire n_3753_o_0;
 wire n_3752_o_0;
 wire n_3751_o_0;
 wire n_3750_o_0;
 wire n_3749_o_0;
 wire n_3748_o_0;
 wire n_3747_o_0;
 wire n_3746_o_0;
 wire n_3745_o_0;
 wire n_3744_o_0;
 wire n_3743_o_0;
 wire n_3742_o_0;
 wire n_3741_o_0;
 wire n_3740_o_0;
 wire n_3739_o_0;
 wire n_3738_o_0;
 wire n_3737_o_0;
 wire n_3736_o_0;
 wire n_3735_o_0;
 wire n_3734_o_0;
 wire n_3733_o_0;
 wire n_3732_o_0;
 wire n_3731_o_0;
 wire n_3730_o_0;
 wire n_3729_o_0;
 wire n_3728_o_0;
 wire n_3727_o_0;
 wire n_3726_o_0;
 wire n_3725_o_0;
 wire n_3724_o_0;
 wire n_3723_o_0;
 wire n_3722_o_0;
 wire n_3721_o_0;
 wire n_3720_o_0;
 wire n_3719_o_0;
 wire n_3718_o_0;
 wire n_3717_o_0;
 wire n_3716_o_0;
 wire n_3715_o_0;
 wire n_3714_o_0;
 wire n_3713_o_0;
 wire n_3712_o_0;
 wire n_3711_o_0;
 wire n_3710_o_0;
 wire n_3709_o_0;
 wire n_3708_o_0;
 wire n_3707_o_0;
 wire n_3706_o_0;
 wire n_3705_o_0;
 wire n_3704_o_0;
 wire n_3703_o_0;
 wire n_3702_o_0;
 wire n_3701_o_0;
 wire n_3700_o_0;
 wire n_3699_o_0;
 wire n_3698_o_0;
 wire n_3697_o_0;
 wire n_3696_o_0;
 wire n_3695_o_0;
 wire n_3694_o_0;
 wire n_3693_o_0;
 wire n_3692_o_0;
 wire n_3691_o_0;
 wire n_3690_o_0;
 wire n_3689_o_0;
 wire n_3688_o_0;
 wire n_3687_o_0;
 wire n_3686_o_0;
 wire n_3685_o_0;
 wire n_3684_o_0;
 wire n_3683_o_0;
 wire n_3682_o_0;
 wire n_3681_o_0;
 wire n_3680_o_0;
 wire n_3679_o_0;
 wire n_3678_o_0;
 wire n_3677_o_0;
 wire n_3676_o_0;
 wire n_3675_o_0;
 wire n_3674_o_0;
 wire n_3673_o_0;
 wire n_3672_o_0;
 wire n_3671_o_0;
 wire n_3670_o_0;
 wire n_3669_o_0;
 wire n_3668_o_0;
 wire n_3667_o_0;
 wire n_3666_o_0;
 wire n_3665_o_0;
 wire n_3664_o_0;
 wire n_3663_o_0;
 wire n_3662_o_0;
 wire n_3661_o_0;
 wire n_3660_o_0;
 wire n_3659_o_0;
 wire n_3658_o_0;
 wire n_3657_o_0;
 wire n_3656_o_0;
 wire n_3655_o_0;
 wire n_3654_o_0;
 wire n_3653_o_0;
 wire n_3652_o_0;
 wire n_3651_o_0;
 wire n_3650_o_0;
 wire n_3649_o_0;
 wire n_3648_o_0;
 wire n_3647_o_0;
 wire n_3646_o_0;
 wire n_3645_o_0;
 wire n_3644_o_0;
 wire n_3643_o_0;
 wire n_3642_o_0;
 wire n_3641_o_0;
 wire n_3640_o_0;
 wire n_3639_o_0;
 wire n_3638_o_0;
 wire n_3637_o_0;
 wire n_3636_o_0;
 wire n_3635_o_0;
 wire n_3634_o_0;
 wire n_3633_o_0;
 wire n_3632_o_0;
 wire n_3631_o_0;
 wire n_3630_o_0;
 wire n_3629_o_0;
 wire n_3628_o_0;
 wire n_3627_o_0;
 wire n_3626_o_0;
 wire n_3625_o_0;
 wire n_3624_o_0;
 wire n_3623_o_0;
 wire n_3622_o_0;
 wire n_3621_o_0;
 wire n_3620_o_0;
 wire n_3619_o_0;
 wire n_3618_o_0;
 wire n_3617_o_0;
 wire n_3616_o_0;
 wire n_3615_o_0;
 wire n_3614_o_0;
 wire n_3613_o_0;
 wire n_3612_o_0;
 wire n_3611_o_0;
 wire n_3610_o_0;
 wire n_3609_o_0;
 wire n_3608_o_0;
 wire n_3607_o_0;
 wire n_3606_o_0;
 wire n_3605_o_0;
 wire n_3604_o_0;
 wire n_3603_o_0;
 wire n_3602_o_0;
 wire n_3601_o_0;
 wire n_3600_o_0;
 wire n_3599_o_0;
 wire n_3598_o_0;
 wire n_3597_o_0;
 wire n_3596_o_0;
 wire n_3595_o_0;
 wire n_3594_o_0;
 wire n_3593_o_0;
 wire n_3592_o_0;
 wire n_3591_o_0;
 wire n_3590_o_0;
 wire n_3589_o_0;
 wire n_3588_o_0;
 wire n_3587_o_0;
 wire n_3586_o_0;
 wire n_3585_o_0;
 wire n_3584_o_0;
 wire n_3583_o_0;
 wire n_3582_o_0;
 wire n_3581_o_0;
 wire n_3580_o_0;
 wire n_3579_o_0;
 wire n_3578_o_0;
 wire n_3577_o_0;
 wire n_3576_o_0;
 wire n_3575_o_0;
 wire n_3574_o_0;
 wire n_3573_o_0;
 wire n_3572_o_0;
 wire n_3571_o_0;
 wire n_3570_o_0;
 wire n_3569_o_0;
 wire n_3568_o_0;
 wire n_3567_o_0;
 wire n_3566_o_0;
 wire n_3565_o_0;
 wire n_3564_o_0;
 wire n_3563_o_0;
 wire n_3562_o_0;
 wire n_3561_o_0;
 wire n_3560_o_0;
 wire n_3559_o_0;
 wire n_3558_o_0;
 wire n_3557_o_0;
 wire n_3556_o_0;
 wire n_3555_o_0;
 wire n_3554_o_0;
 wire n_3553_o_0;
 wire n_3552_o_0;
 wire n_3551_o_0;
 wire n_3550_o_0;
 wire n_3549_o_0;
 wire n_3548_o_0;
 wire n_3547_o_0;
 wire n_3546_o_0;
 wire n_3545_o_0;
 wire n_3544_o_0;
 wire n_3543_o_0;
 wire n_3542_o_0;
 wire n_3541_o_0;
 wire n_3540_o_0;
 wire n_3539_o_0;
 wire n_3538_o_0;
 wire n_3537_o_0;
 wire n_3536_o_0;
 wire n_3535_o_0;
 wire n_3534_o_0;
 wire n_3533_o_0;
 wire n_3532_o_0;
 wire n_3531_o_0;
 wire n_3530_o_0;
 wire n_3529_o_0;
 wire n_3528_o_0;
 wire n_3527_o_0;
 wire n_3526_o_0;
 wire n_3525_o_0;
 wire n_3524_o_0;
 wire n_3523_o_0;
 wire n_3522_o_0;
 wire n_3521_o_0;
 wire n_3520_o_0;
 wire n_3519_o_0;
 wire n_3518_o_0;
 wire n_3517_o_0;
 wire n_3516_o_0;
 wire n_3515_o_0;
 wire n_3514_o_0;
 wire n_3513_o_0;
 wire n_3512_o_0;
 wire n_3511_o_0;
 wire n_3510_o_0;
 wire n_3509_o_0;
 wire n_3508_o_0;
 wire n_3507_o_0;
 wire n_3506_o_0;
 wire n_3505_o_0;
 wire n_3504_o_0;
 wire n_3503_o_0;
 wire n_3502_o_0;
 wire n_3501_o_0;
 wire n_3500_o_0;
 wire n_3499_o_0;
 wire n_3498_o_0;
 wire n_3497_o_0;
 wire n_3496_o_0;
 wire n_3495_o_0;
 wire n_3494_o_0;
 wire n_3493_o_0;
 wire n_3492_o_0;
 wire n_3491_o_0;
 wire n_3490_o_0;
 wire n_3489_o_0;
 wire n_3488_o_0;
 wire n_3487_o_0;
 wire n_3486_o_0;
 wire n_3485_o_0;
 wire n_3484_o_0;
 wire n_3483_o_0;
 wire n_3482_o_0;
 wire n_3481_o_0;
 wire n_3480_o_0;
 wire n_3479_o_0;
 wire n_3478_o_0;
 wire n_3477_o_0;
 wire n_3476_o_0;
 wire n_3475_o_0;
 wire n_3474_o_0;
 wire n_3473_o_0;
 wire n_3472_o_0;
 wire n_3471_o_0;
 wire n_3470_o_0;
 wire n_3469_o_0;
 wire n_3468_o_0;
 wire n_3467_o_0;
 wire n_3466_o_0;
 wire n_3465_o_0;
 wire n_3464_o_0;
 wire n_3463_o_0;
 wire n_3462_o_0;
 wire n_3461_o_0;
 wire n_3460_o_0;
 wire n_3459_o_0;
 wire n_3458_o_0;
 wire n_3457_o_0;
 wire n_3456_o_0;
 wire n_3455_o_0;
 wire n_3454_o_0;
 wire n_3453_o_0;
 wire n_3452_o_0;
 wire n_3451_o_0;
 wire n_3450_o_0;
 wire n_3449_o_0;
 wire n_3448_o_0;
 wire n_3447_o_0;
 wire n_3446_o_0;
 wire n_3445_o_0;
 wire n_3444_o_0;
 wire n_3443_o_0;
 wire n_3442_o_0;
 wire n_3441_o_0;
 wire n_3440_o_0;
 wire n_3439_o_0;
 wire n_3438_o_0;
 wire n_3437_o_0;
 wire n_3436_o_0;
 wire n_3435_o_0;
 wire n_3434_o_0;
 wire n_3433_o_0;
 wire n_3432_o_0;
 wire n_3431_o_0;
 wire n_3430_o_0;
 wire n_3429_o_0;
 wire n_3428_o_0;
 wire n_3427_o_0;
 wire n_3426_o_0;
 wire n_3425_o_0;
 wire n_3424_o_0;
 wire n_3423_o_0;
 wire n_3422_o_0;
 wire n_3421_o_0;
 wire n_3420_o_0;
 wire n_3419_o_0;
 wire n_3418_o_0;
 wire n_3417_o_0;
 wire n_3416_o_0;
 wire n_3415_o_0;
 wire n_3414_o_0;
 wire n_3413_o_0;
 wire n_3412_o_0;
 wire n_3411_o_0;
 wire n_3410_o_0;
 wire n_3409_o_0;
 wire n_3408_o_0;
 wire n_3407_o_0;
 wire n_3406_o_0;
 wire n_3405_o_0;
 wire n_3404_o_0;
 wire n_3403_o_0;
 wire n_3402_o_0;
 wire n_3401_o_0;
 wire n_3400_o_0;
 wire n_3399_o_0;
 wire n_3398_o_0;
 wire n_3397_o_0;
 wire n_3396_o_0;
 wire n_3395_o_0;
 wire n_3394_o_0;
 wire n_3393_o_0;
 wire n_3392_o_0;
 wire n_3391_o_0;
 wire n_3390_o_0;
 wire n_3389_o_0;
 wire n_3388_o_0;
 wire n_3387_o_0;
 wire n_3386_o_0;
 wire n_3385_o_0;
 wire n_3384_o_0;
 wire n_3383_o_0;
 wire n_3382_o_0;
 wire n_3381_o_0;
 wire n_3380_o_0;
 wire n_3379_o_0;
 wire n_3378_o_0;
 wire n_3377_o_0;
 wire n_3376_o_0;
 wire n_3375_o_0;
 wire n_3374_o_0;
 wire n_3373_o_0;
 wire n_3372_o_0;
 wire n_3371_o_0;
 wire n_3370_o_0;
 wire n_3369_o_0;
 wire n_3368_o_0;
 wire n_3367_o_0;
 wire n_3366_o_0;
 wire n_3365_o_0;
 wire n_3364_o_0;
 wire n_3363_o_0;
 wire n_3362_o_0;
 wire n_3361_o_0;
 wire n_3360_o_0;
 wire n_3359_o_0;
 wire n_3358_o_0;
 wire n_3357_o_0;
 wire n_3356_o_0;
 wire n_3355_o_0;
 wire n_3354_o_0;
 wire n_3353_o_0;
 wire n_3352_o_0;
 wire n_3351_o_0;
 wire n_3350_o_0;
 wire n_3349_o_0;
 wire n_3348_o_0;
 wire n_3347_o_0;
 wire n_3346_o_0;
 wire n_3345_o_0;
 wire n_3344_o_0;
 wire n_3343_o_0;
 wire n_3342_o_0;
 wire n_3341_o_0;
 wire n_3340_o_0;
 wire n_3339_o_0;
 wire n_3338_o_0;
 wire n_3337_o_0;
 wire n_3336_o_0;
 wire n_3335_o_0;
 wire n_3334_o_0;
 wire n_3333_o_0;
 wire n_3332_o_0;
 wire n_3331_o_0;
 wire n_3330_o_0;
 wire n_3329_o_0;
 wire n_3328_o_0;
 wire n_3327_o_0;
 wire n_3326_o_0;
 wire n_3325_o_0;
 wire n_3324_o_0;
 wire n_3323_o_0;
 wire n_3322_o_0;
 wire n_3321_o_0;
 wire n_3320_o_0;
 wire n_3319_o_0;
 wire n_3318_o_0;
 wire n_3317_o_0;
 wire n_3316_o_0;
 wire n_3315_o_0;
 wire n_3314_o_0;
 wire n_3313_o_0;
 wire n_3312_o_0;
 wire n_3311_o_0;
 wire n_3310_o_0;
 wire n_3309_o_0;
 wire n_3308_o_0;
 wire n_3307_o_0;
 wire n_3306_o_0;
 wire n_3305_o_0;
 wire n_3304_o_0;
 wire n_3303_o_0;
 wire n_3302_o_0;
 wire n_3301_o_0;
 wire n_3300_o_0;
 wire n_3299_o_0;
 wire n_3298_o_0;
 wire n_3297_o_0;
 wire n_3296_o_0;
 wire n_3295_o_0;
 wire n_3294_o_0;
 wire n_3293_o_0;
 wire n_3292_o_0;
 wire n_3291_o_0;
 wire n_3290_o_0;
 wire n_3289_o_0;
 wire n_3288_o_0;
 wire n_3287_o_0;
 wire n_3286_o_0;
 wire n_3285_o_0;
 wire n_3284_o_0;
 wire n_3283_o_0;
 wire n_3282_o_0;
 wire n_3281_o_0;
 wire n_3280_o_0;
 wire n_3279_o_0;
 wire n_3278_o_0;
 wire n_3277_o_0;
 wire n_3276_o_0;
 wire n_3275_o_0;
 wire n_3274_o_0;
 wire n_3273_o_0;
 wire n_3272_o_0;
 wire n_3271_o_0;
 wire n_3270_o_0;
 wire n_3269_o_0;
 wire n_3268_o_0;
 wire n_3267_o_0;
 wire n_3266_o_0;
 wire n_3265_o_0;
 wire n_3264_o_0;
 wire n_3263_o_0;
 wire n_3262_o_0;
 wire n_3261_o_0;
 wire n_3260_o_0;
 wire n_3259_o_0;
 wire n_3258_o_0;
 wire n_3257_o_0;
 wire n_3256_o_0;
 wire n_3255_o_0;
 wire n_3254_o_0;
 wire n_3253_o_0;
 wire n_3252_o_0;
 wire n_3251_o_0;
 wire n_3250_o_0;
 wire n_3249_o_0;
 wire n_3248_o_0;
 wire n_3247_o_0;
 wire n_3246_o_0;
 wire n_3245_o_0;
 wire n_3244_o_0;
 wire n_3243_o_0;
 wire n_3242_o_0;
 wire n_3241_o_0;
 wire n_3240_o_0;
 wire n_3239_o_0;
 wire n_3238_o_0;
 wire n_3237_o_0;
 wire n_3236_o_0;
 wire n_3235_o_0;
 wire n_3234_o_0;
 wire n_3233_o_0;
 wire n_3232_o_0;
 wire n_3231_o_0;
 wire n_3230_o_0;
 wire n_3229_o_0;
 wire n_3228_o_0;
 wire n_3227_o_0;
 wire n_3226_o_0;
 wire n_3225_o_0;
 wire n_3224_o_0;
 wire n_3223_o_0;
 wire n_3222_o_0;
 wire n_3221_o_0;
 wire n_3220_o_0;
 wire n_3219_o_0;
 wire n_3218_o_0;
 wire n_3217_o_0;
 wire n_3216_o_0;
 wire n_3215_o_0;
 wire n_3214_o_0;
 wire n_3213_o_0;
 wire n_3212_o_0;
 wire n_3211_o_0;
 wire n_3210_o_0;
 wire n_3209_o_0;
 wire n_3208_o_0;
 wire n_3207_o_0;
 wire n_3206_o_0;
 wire n_3205_o_0;
 wire n_3204_o_0;
 wire n_3203_o_0;
 wire n_3202_o_0;
 wire n_3201_o_0;
 wire n_3200_o_0;
 wire n_3199_o_0;
 wire n_3198_o_0;
 wire n_3197_o_0;
 wire n_3196_o_0;
 wire n_3195_o_0;
 wire n_3194_o_0;
 wire n_3193_o_0;
 wire n_3192_o_0;
 wire n_3191_o_0;
 wire n_3190_o_0;
 wire n_3189_o_0;
 wire n_3188_o_0;
 wire n_3187_o_0;
 wire n_3186_o_0;
 wire n_3185_o_0;
 wire n_3184_o_0;
 wire n_3183_o_0;
 wire n_3182_o_0;
 wire n_3181_o_0;
 wire n_3180_o_0;
 wire n_3179_o_0;
 wire n_3178_o_0;
 wire n_3177_o_0;
 wire n_3176_o_0;
 wire n_3175_o_0;
 wire n_3174_o_0;
 wire n_3173_o_0;
 wire n_3172_o_0;
 wire n_3171_o_0;
 wire n_3170_o_0;
 wire n_3169_o_0;
 wire n_3168_o_0;
 wire n_3167_o_0;
 wire n_3166_o_0;
 wire n_3165_o_0;
 wire n_3164_o_0;
 wire n_3163_o_0;
 wire n_3162_o_0;
 wire n_3161_o_0;
 wire n_3160_o_0;
 wire n_3159_o_0;
 wire n_3158_o_0;
 wire n_3157_o_0;
 wire n_3156_o_0;
 wire n_3155_o_0;
 wire n_3154_o_0;
 wire n_3153_o_0;
 wire n_3152_o_0;
 wire n_3151_o_0;
 wire n_3150_o_0;
 wire n_3149_o_0;
 wire n_3148_o_0;
 wire n_3147_o_0;
 wire n_3146_o_0;
 wire n_3145_o_0;
 wire n_3144_o_0;
 wire n_3143_o_0;
 wire n_3142_o_0;
 wire n_3141_o_0;
 wire n_3140_o_0;
 wire n_3139_o_0;
 wire n_3138_o_0;
 wire n_3137_o_0;
 wire n_3136_o_0;
 wire n_3135_o_0;
 wire n_3134_o_0;
 wire n_3133_o_0;
 wire n_3132_o_0;
 wire n_3131_o_0;
 wire n_3130_o_0;
 wire n_3129_o_0;
 wire n_3128_o_0;
 wire n_3127_o_0;
 wire n_3126_o_0;
 wire n_3125_o_0;
 wire n_3124_o_0;
 wire n_3123_o_0;
 wire n_3122_o_0;
 wire n_3121_o_0;
 wire n_3120_o_0;
 wire n_3119_o_0;
 wire n_3118_o_0;
 wire n_3117_o_0;
 wire n_3116_o_0;
 wire n_3115_o_0;
 wire n_3114_o_0;
 wire n_3113_o_0;
 wire n_3112_o_0;
 wire n_3111_o_0;
 wire n_3110_o_0;
 wire n_3109_o_0;
 wire n_3108_o_0;
 wire n_3107_o_0;
 wire n_3106_o_0;
 wire n_3105_o_0;
 wire n_3104_o_0;
 wire n_3103_o_0;
 wire n_3102_o_0;
 wire n_3101_o_0;
 wire n_3100_o_0;
 wire n_3099_o_0;
 wire n_3098_o_0;
 wire n_3097_o_0;
 wire n_3096_o_0;
 wire n_3095_o_0;
 wire n_3094_o_0;
 wire n_3093_o_0;
 wire n_3092_o_0;
 wire n_3091_o_0;
 wire n_3090_o_0;
 wire n_3089_o_0;
 wire n_3088_o_0;
 wire n_3087_o_0;
 wire n_3086_o_0;
 wire n_3085_o_0;
 wire n_3084_o_0;
 wire n_3083_o_0;
 wire n_3082_o_0;
 wire n_3081_o_0;
 wire n_3080_o_0;
 wire n_3079_o_0;
 wire n_3078_o_0;
 wire n_3077_o_0;
 wire n_3076_o_0;
 wire n_3075_o_0;
 wire n_3074_o_0;
 wire n_3073_o_0;
 wire n_3072_o_0;
 wire n_3071_o_0;
 wire n_3070_o_0;
 wire n_3069_o_0;
 wire n_3068_o_0;
 wire n_3067_o_0;
 wire n_3066_o_0;
 wire n_3065_o_0;
 wire n_3064_o_0;
 wire n_3063_o_0;
 wire n_3062_o_0;
 wire n_3061_o_0;
 wire n_3060_o_0;
 wire n_3059_o_0;
 wire n_3058_o_0;
 wire n_3057_o_0;
 wire n_3056_o_0;
 wire n_3055_o_0;
 wire n_3054_o_0;
 wire n_3053_o_0;
 wire n_3052_o_0;
 wire n_3051_o_0;
 wire n_3050_o_0;
 wire n_3049_o_0;
 wire n_3048_o_0;
 wire n_3047_o_0;
 wire n_3046_o_0;
 wire n_3045_o_0;
 wire n_3044_o_0;
 wire n_3043_o_0;
 wire n_3042_o_0;
 wire n_3041_o_0;
 wire n_3040_o_0;
 wire n_3039_o_0;
 wire n_3038_o_0;
 wire n_3037_o_0;
 wire n_3036_o_0;
 wire n_3035_o_0;
 wire n_3034_o_0;
 wire n_3033_o_0;
 wire n_3032_o_0;
 wire n_3031_o_0;
 wire n_3030_o_0;
 wire n_3029_o_0;
 wire n_3028_o_0;
 wire n_3027_o_0;
 wire n_3026_o_0;
 wire n_3025_o_0;
 wire n_3024_o_0;
 wire n_3023_o_0;
 wire n_3022_o_0;
 wire n_3021_o_0;
 wire n_3020_o_0;
 wire n_3019_o_0;
 wire n_3018_o_0;
 wire n_3017_o_0;
 wire n_3016_o_0;
 wire n_3015_o_0;
 wire n_3014_o_0;
 wire n_3013_o_0;
 wire n_3012_o_0;
 wire n_3011_o_0;
 wire n_3010_o_0;
 wire n_3009_o_0;
 wire n_3008_o_0;
 wire n_3007_o_0;
 wire n_3006_o_0;
 wire n_3005_o_0;
 wire n_3004_o_0;
 wire n_3003_o_0;
 wire n_3002_o_0;
 wire n_3001_o_0;
 wire n_3000_o_0;
 wire n_2999_o_0;
 wire n_2998_o_0;
 wire n_2997_o_0;
 wire n_2996_o_0;
 wire n_2995_o_0;
 wire n_2994_o_0;
 wire n_2993_o_0;
 wire n_2992_o_0;
 wire n_2991_o_0;
 wire n_2990_o_0;
 wire n_2989_o_0;
 wire n_2988_o_0;
 wire n_2987_o_0;
 wire n_2986_o_0;
 wire n_2985_o_0;
 wire n_2984_o_0;
 wire n_2983_o_0;
 wire n_2982_o_0;
 wire n_2981_o_0;
 wire n_2980_o_0;
 wire n_2979_o_0;
 wire n_2978_o_0;
 wire n_2977_o_0;
 wire n_2976_o_0;
 wire n_2975_o_0;
 wire n_2974_o_0;
 wire n_2973_o_0;
 wire n_2972_o_0;
 wire n_2971_o_0;
 wire n_2970_o_0;
 wire n_2969_o_0;
 wire n_2968_o_0;
 wire n_2967_o_0;
 wire n_2966_o_0;
 wire n_2965_o_0;
 wire n_2964_o_0;
 wire n_2963_o_0;
 wire n_2962_o_0;
 wire n_2961_o_0;
 wire n_2960_o_0;
 wire n_2959_o_0;
 wire n_2958_o_0;
 wire n_2957_o_0;
 wire n_2956_o_0;
 wire n_2955_o_0;
 wire n_2954_o_0;
 wire n_2953_o_0;
 wire n_2952_o_0;
 wire n_2951_o_0;
 wire n_2950_o_0;
 wire n_2949_o_0;
 wire n_2948_o_0;
 wire n_2947_o_0;
 wire n_2946_o_0;
 wire n_2945_o_0;
 wire n_2944_o_0;
 wire n_2943_o_0;
 wire n_2942_o_0;
 wire n_2941_o_0;
 wire n_2940_o_0;
 wire n_2939_o_0;
 wire n_2938_o_0;
 wire n_2937_o_0;
 wire n_2936_o_0;
 wire n_2935_o_0;
 wire n_2934_o_0;
 wire n_2933_o_0;
 wire n_2932_o_0;
 wire n_2931_o_0;
 wire n_2930_o_0;
 wire n_2929_o_0;
 wire n_2928_o_0;
 wire n_2927_o_0;
 wire n_2926_o_0;
 wire n_2925_o_0;
 wire n_2924_o_0;
 wire n_2923_o_0;
 wire n_2922_o_0;
 wire n_2921_o_0;
 wire n_2920_o_0;
 wire n_2919_o_0;
 wire n_2918_o_0;
 wire n_2917_o_0;
 wire n_2916_o_0;
 wire n_2915_o_0;
 wire n_2914_o_0;
 wire n_2913_o_0;
 wire n_2912_o_0;
 wire n_2911_o_0;
 wire n_2910_o_0;
 wire n_2909_o_0;
 wire n_2908_o_0;
 wire n_2907_o_0;
 wire n_2906_o_0;
 wire n_2905_o_0;
 wire n_2904_o_0;
 wire n_2903_o_0;
 wire n_2902_o_0;
 wire n_2901_o_0;
 wire n_2900_o_0;
 wire n_2899_o_0;
 wire n_2898_o_0;
 wire n_2897_o_0;
 wire n_2896_o_0;
 wire n_2895_o_0;
 wire n_2894_o_0;
 wire n_2893_o_0;
 wire n_2892_o_0;
 wire n_2891_o_0;
 wire n_2890_o_0;
 wire n_2889_o_0;
 wire n_2888_o_0;
 wire n_2887_o_0;
 wire n_2886_o_0;
 wire n_2885_o_0;
 wire n_2884_o_0;
 wire n_2883_o_0;
 wire n_2882_o_0;
 wire n_2881_o_0;
 wire n_2880_o_0;
 wire n_2879_o_0;
 wire n_2878_o_0;
 wire n_2877_o_0;
 wire n_2876_o_0;
 wire n_2875_o_0;
 wire n_2874_o_0;
 wire n_2873_o_0;
 wire n_2872_o_0;
 wire n_2871_o_0;
 wire n_2870_o_0;
 wire n_2869_o_0;
 wire n_2868_o_0;
 wire n_2867_o_0;
 wire n_2866_o_0;
 wire n_2865_o_0;
 wire n_2864_o_0;
 wire n_2863_o_0;
 wire n_2862_o_0;
 wire n_2861_o_0;
 wire n_2860_o_0;
 wire n_2859_o_0;
 wire n_2858_o_0;
 wire n_2857_o_0;
 wire n_2856_o_0;
 wire n_2855_o_0;
 wire n_2854_o_0;
 wire n_2853_o_0;
 wire n_2852_o_0;
 wire n_2851_o_0;
 wire n_2850_o_0;
 wire n_2849_o_0;
 wire n_2848_o_0;
 wire n_2847_o_0;
 wire n_2846_o_0;
 wire n_2845_o_0;
 wire n_2844_o_0;
 wire n_2843_o_0;
 wire n_2842_o_0;
 wire n_2841_o_0;
 wire n_2840_o_0;
 wire n_2839_o_0;
 wire n_2838_o_0;
 wire n_2837_o_0;
 wire n_2836_o_0;
 wire n_2835_o_0;
 wire n_2834_o_0;
 wire n_2833_o_0;
 wire n_2832_o_0;
 wire n_2831_o_0;
 wire n_2830_o_0;
 wire n_2829_o_0;
 wire n_2828_o_0;
 wire n_2827_o_0;
 wire n_2826_o_0;
 wire n_2825_o_0;
 wire n_2824_o_0;
 wire n_2823_o_0;
 wire n_2822_o_0;
 wire n_2821_o_0;
 wire n_2820_o_0;
 wire n_2819_o_0;
 wire n_2818_o_0;
 wire n_2817_o_0;
 wire n_2816_o_0;
 wire n_2815_o_0;
 wire n_2814_o_0;
 wire n_2813_o_0;
 wire n_2812_o_0;
 wire n_2811_o_0;
 wire n_2810_o_0;
 wire n_2809_o_0;
 wire n_2808_o_0;
 wire n_2807_o_0;
 wire n_2806_o_0;
 wire n_2805_o_0;
 wire n_2804_o_0;
 wire n_2803_o_0;
 wire n_2802_o_0;
 wire n_2801_o_0;
 wire n_2800_o_0;
 wire n_2799_o_0;
 wire n_2798_o_0;
 wire n_2797_o_0;
 wire n_2796_o_0;
 wire n_2795_o_0;
 wire n_2794_o_0;
 wire n_2793_o_0;
 wire n_2792_o_0;
 wire n_2791_o_0;
 wire n_2790_o_0;
 wire n_2789_o_0;
 wire n_2788_o_0;
 wire n_2787_o_0;
 wire n_2786_o_0;
 wire n_2785_o_0;
 wire n_2784_o_0;
 wire n_2783_o_0;
 wire n_2782_o_0;
 wire n_2781_o_0;
 wire n_2780_o_0;
 wire n_2779_o_0;
 wire n_2778_o_0;
 wire n_2777_o_0;
 wire n_2776_o_0;
 wire n_2775_o_0;
 wire n_2774_o_0;
 wire n_2773_o_0;
 wire n_2772_o_0;
 wire n_2771_o_0;
 wire n_2770_o_0;
 wire n_2769_o_0;
 wire n_2768_o_0;
 wire n_2767_o_0;
 wire n_2766_o_0;
 wire n_2765_o_0;
 wire n_2764_o_0;
 wire n_2763_o_0;
 wire n_2762_o_0;
 wire n_2761_o_0;
 wire n_2760_o_0;
 wire n_2759_o_0;
 wire n_2758_o_0;
 wire n_2757_o_0;
 wire n_2756_o_0;
 wire n_2755_o_0;
 wire n_2754_o_0;
 wire n_2753_o_0;
 wire n_2752_o_0;
 wire n_2751_o_0;
 wire n_2750_o_0;
 wire n_2749_o_0;
 wire n_2748_o_0;
 wire n_2747_o_0;
 wire n_2746_o_0;
 wire n_2745_o_0;
 wire n_2744_o_0;
 wire n_2743_o_0;
 wire n_2742_o_0;
 wire n_2741_o_0;
 wire n_2740_o_0;
 wire n_2739_o_0;
 wire n_2738_o_0;
 wire n_2737_o_0;
 wire n_2736_o_0;
 wire n_2735_o_0;
 wire n_2734_o_0;
 wire n_2733_o_0;
 wire n_2732_o_0;
 wire n_2731_o_0;
 wire n_2730_o_0;
 wire n_2729_o_0;
 wire n_2728_o_0;
 wire n_2727_o_0;
 wire n_2726_o_0;
 wire n_2725_o_0;
 wire n_2724_o_0;
 wire n_2723_o_0;
 wire n_2722_o_0;
 wire n_2721_o_0;
 wire n_2720_o_0;
 wire n_2719_o_0;
 wire n_2718_o_0;
 wire n_2717_o_0;
 wire n_2716_o_0;
 wire n_2715_o_0;
 wire n_2714_o_0;
 wire n_2713_o_0;
 wire n_2712_o_0;
 wire n_2711_o_0;
 wire n_2710_o_0;
 wire n_2709_o_0;
 wire n_2708_o_0;
 wire n_2707_o_0;
 wire n_2706_o_0;
 wire n_2705_o_0;
 wire n_2704_o_0;
 wire n_2703_o_0;
 wire n_2702_o_0;
 wire n_2701_o_0;
 wire n_2700_o_0;
 wire n_2699_o_0;
 wire n_2698_o_0;
 wire n_2697_o_0;
 wire n_2696_o_0;
 wire n_2695_o_0;
 wire n_2694_o_0;
 wire n_2693_o_0;
 wire n_2692_o_0;
 wire n_2691_o_0;
 wire n_2690_o_0;
 wire n_2689_o_0;
 wire n_2688_o_0;
 wire n_2687_o_0;
 wire n_2686_o_0;
 wire n_2685_o_0;
 wire n_2684_o_0;
 wire n_2683_o_0;
 wire n_2682_o_0;
 wire n_2681_o_0;
 wire n_2680_o_0;
 wire n_2679_o_0;
 wire n_2678_o_0;
 wire n_2677_o_0;
 wire n_2676_o_0;
 wire n_2675_o_0;
 wire n_2674_o_0;
 wire n_2673_o_0;
 wire n_2672_o_0;
 wire n_2671_o_0;
 wire n_2670_o_0;
 wire n_2669_o_0;
 wire n_2668_o_0;
 wire n_2667_o_0;
 wire n_2666_o_0;
 wire n_2665_o_0;
 wire n_2664_o_0;
 wire n_2663_o_0;
 wire n_2662_o_0;
 wire n_2661_o_0;
 wire n_2660_o_0;
 wire n_2659_o_0;
 wire n_2658_o_0;
 wire n_2657_o_0;
 wire n_2656_o_0;
 wire n_2655_o_0;
 wire n_2654_o_0;
 wire n_2653_o_0;
 wire n_2652_o_0;
 wire n_2651_o_0;
 wire n_2650_o_0;
 wire n_2649_o_0;
 wire n_2648_o_0;
 wire n_2647_o_0;
 wire n_2646_o_0;
 wire n_2645_o_0;
 wire n_2644_o_0;
 wire n_2643_o_0;
 wire n_2642_o_0;
 wire n_2641_o_0;
 wire n_2640_o_0;
 wire n_2639_o_0;
 wire n_2638_o_0;
 wire n_2637_o_0;
 wire n_2636_o_0;
 wire n_2635_o_0;
 wire n_2634_o_0;
 wire n_2633_o_0;
 wire n_2632_o_0;
 wire n_2631_o_0;
 wire n_2630_o_0;
 wire n_2629_o_0;
 wire n_2628_o_0;
 wire n_2627_o_0;
 wire n_2626_o_0;
 wire n_2625_o_0;
 wire n_2624_o_0;
 wire n_2623_o_0;
 wire n_2622_o_0;
 wire n_2621_o_0;
 wire n_2620_o_0;
 wire n_2619_o_0;
 wire n_2618_o_0;
 wire n_2617_o_0;
 wire n_2616_o_0;
 wire n_2615_o_0;
 wire n_2614_o_0;
 wire n_2613_o_0;
 wire n_2612_o_0;
 wire n_2611_o_0;
 wire n_2610_o_0;
 wire n_2609_o_0;
 wire n_2608_o_0;
 wire n_2607_o_0;
 wire n_2606_o_0;
 wire n_2605_o_0;
 wire n_2604_o_0;
 wire n_2603_o_0;
 wire n_2602_o_0;
 wire n_2601_o_0;
 wire n_2600_o_0;
 wire n_2599_o_0;
 wire n_2598_o_0;
 wire n_2597_o_0;
 wire n_2596_o_0;
 wire n_2595_o_0;
 wire n_2594_o_0;
 wire n_2593_o_0;
 wire n_2592_o_0;
 wire n_2591_o_0;
 wire n_2590_o_0;
 wire n_2589_o_0;
 wire n_2588_o_0;
 wire n_2587_o_0;
 wire n_2586_o_0;
 wire n_2585_o_0;
 wire n_2584_o_0;
 wire n_2583_o_0;
 wire n_2582_o_0;
 wire n_2581_o_0;
 wire n_2580_o_0;
 wire n_2579_o_0;
 wire n_2578_o_0;
 wire n_2577_o_0;
 wire n_2576_o_0;
 wire n_2575_o_0;
 wire n_2574_o_0;
 wire n_2573_o_0;
 wire n_2572_o_0;
 wire n_2571_o_0;
 wire n_2570_o_0;
 wire n_2569_o_0;
 wire n_2568_o_0;
 wire n_2567_o_0;
 wire n_2566_o_0;
 wire n_2565_o_0;
 wire n_2564_o_0;
 wire n_2563_o_0;
 wire n_2562_o_0;
 wire n_2561_o_0;
 wire n_2560_o_0;
 wire n_2559_o_0;
 wire n_2558_o_0;
 wire n_2557_o_0;
 wire n_2556_o_0;
 wire n_2555_o_0;
 wire n_2554_o_0;
 wire n_2553_o_0;
 wire n_2552_o_0;
 wire n_2551_o_0;
 wire n_2550_o_0;
 wire n_2549_o_0;
 wire n_2548_o_0;
 wire n_2547_o_0;
 wire n_2546_o_0;
 wire n_2545_o_0;
 wire n_2544_o_0;
 wire n_2543_o_0;
 wire n_2542_o_0;
 wire n_2541_o_0;
 wire n_2540_o_0;
 wire n_2539_o_0;
 wire n_2538_o_0;
 wire n_2537_o_0;
 wire n_2536_o_0;
 wire n_2535_o_0;
 wire n_2534_o_0;
 wire n_2533_o_0;
 wire n_2532_o_0;
 wire n_2531_o_0;
 wire n_2530_o_0;
 wire n_2529_o_0;
 wire n_2528_o_0;
 wire n_2527_o_0;
 wire n_2526_o_0;
 wire n_2525_o_0;
 wire n_2524_o_0;
 wire n_2523_o_0;
 wire n_2522_o_0;
 wire n_2521_o_0;
 wire n_2520_o_0;
 wire n_2519_o_0;
 wire n_2518_o_0;
 wire n_2517_o_0;
 wire n_2516_o_0;
 wire n_2515_o_0;
 wire n_2514_o_0;
 wire n_2513_o_0;
 wire n_2512_o_0;
 wire n_2511_o_0;
 wire n_2510_o_0;
 wire n_2509_o_0;
 wire n_2508_o_0;
 wire n_2507_o_0;
 wire n_2506_o_0;
 wire n_2505_o_0;
 wire n_2504_o_0;
 wire n_2503_o_0;
 wire n_2502_o_0;
 wire n_2501_o_0;
 wire n_2500_o_0;
 wire n_2499_o_0;
 wire n_2498_o_0;
 wire n_2497_o_0;
 wire n_2496_o_0;
 wire n_2495_o_0;
 wire n_2494_o_0;
 wire n_2493_o_0;
 wire n_2492_o_0;
 wire n_2491_o_0;
 wire n_2490_o_0;
 wire n_2489_o_0;
 wire n_2488_o_0;
 wire n_2487_o_0;
 wire n_2486_o_0;
 wire n_2485_o_0;
 wire n_2484_o_0;
 wire n_2483_o_0;
 wire n_2482_o_0;
 wire n_2481_o_0;
 wire n_2480_o_0;
 wire n_2479_o_0;
 wire n_2478_o_0;
 wire n_2477_o_0;
 wire n_2476_o_0;
 wire n_2475_o_0;
 wire n_2474_o_0;
 wire n_2473_o_0;
 wire n_2472_o_0;
 wire n_2471_o_0;
 wire n_2470_o_0;
 wire n_2469_o_0;
 wire n_2468_o_0;
 wire n_2467_o_0;
 wire n_2466_o_0;
 wire n_2465_o_0;
 wire n_2464_o_0;
 wire n_2463_o_0;
 wire n_2462_o_0;
 wire n_2461_o_0;
 wire n_2460_o_0;
 wire n_2459_o_0;
 wire n_2458_o_0;
 wire n_2457_o_0;
 wire n_2456_o_0;
 wire n_2455_o_0;
 wire n_2454_o_0;
 wire n_2453_o_0;
 wire n_2452_o_0;
 wire n_2451_o_0;
 wire n_2450_o_0;
 wire n_2449_o_0;
 wire n_2448_o_0;
 wire n_2447_o_0;
 wire n_2446_o_0;
 wire n_2445_o_0;
 wire n_2444_o_0;
 wire n_2443_o_0;
 wire n_2442_o_0;
 wire n_2441_o_0;
 wire n_2440_o_0;
 wire n_2439_o_0;
 wire n_2438_o_0;
 wire n_2437_o_0;
 wire n_2436_o_0;
 wire n_2435_o_0;
 wire n_2434_o_0;
 wire n_2433_o_0;
 wire n_2432_o_0;
 wire n_2431_o_0;
 wire n_2430_o_0;
 wire n_2429_o_0;
 wire n_2428_o_0;
 wire n_2427_o_0;
 wire n_2426_o_0;
 wire n_2425_o_0;
 wire n_2424_o_0;
 wire n_2423_o_0;
 wire n_2422_o_0;
 wire n_2421_o_0;
 wire n_2420_o_0;
 wire n_2419_o_0;
 wire n_2418_o_0;
 wire n_2417_o_0;
 wire n_2416_o_0;
 wire n_2415_o_0;
 wire n_2414_o_0;
 wire n_2413_o_0;
 wire n_2412_o_0;
 wire n_2411_o_0;
 wire n_2410_o_0;
 wire n_2409_o_0;
 wire n_2408_o_0;
 wire n_2407_o_0;
 wire n_2406_o_0;
 wire n_2405_o_0;
 wire n_2404_o_0;
 wire n_2403_o_0;
 wire n_2402_o_0;
 wire n_2401_o_0;
 wire n_2400_o_0;
 wire n_2399_o_0;
 wire n_2398_o_0;
 wire n_2397_o_0;
 wire n_2396_o_0;
 wire n_2395_o_0;
 wire n_2394_o_0;
 wire n_2393_o_0;
 wire n_2392_o_0;
 wire n_2391_o_0;
 wire n_2390_o_0;
 wire n_2389_o_0;
 wire n_2388_o_0;
 wire n_2387_o_0;
 wire n_2386_o_0;
 wire n_2385_o_0;
 wire n_2384_o_0;
 wire n_2383_o_0;
 wire n_2382_o_0;
 wire n_2381_o_0;
 wire n_2380_o_0;
 wire n_2379_o_0;
 wire n_2378_o_0;
 wire n_2377_o_0;
 wire n_2376_o_0;
 wire n_2375_o_0;
 wire n_2374_o_0;
 wire n_2373_o_0;
 wire n_2372_o_0;
 wire n_2371_o_0;
 wire n_2370_o_0;
 wire n_2369_o_0;
 wire n_2368_o_0;
 wire n_2367_o_0;
 wire n_2366_o_0;
 wire n_2365_o_0;
 wire n_2364_o_0;
 wire n_2363_o_0;
 wire n_2362_o_0;
 wire n_2361_o_0;
 wire n_2360_o_0;
 wire n_2359_o_0;
 wire n_2358_o_0;
 wire n_2357_o_0;
 wire n_2356_o_0;
 wire n_2355_o_0;
 wire n_2354_o_0;
 wire n_2353_o_0;
 wire n_2352_o_0;
 wire n_2351_o_0;
 wire n_2350_o_0;
 wire n_2349_o_0;
 wire n_2348_o_0;
 wire n_2347_o_0;
 wire n_2346_o_0;
 wire n_2345_o_0;
 wire n_2344_o_0;
 wire n_2343_o_0;
 wire n_2342_o_0;
 wire n_2341_o_0;
 wire n_2340_o_0;
 wire n_2339_o_0;
 wire n_2338_o_0;
 wire n_2337_o_0;
 wire n_2336_o_0;
 wire n_2335_o_0;
 wire n_2334_o_0;
 wire n_2333_o_0;
 wire n_2332_o_0;
 wire n_2331_o_0;
 wire n_2330_o_0;
 wire n_2329_o_0;
 wire n_2328_o_0;
 wire n_2327_o_0;
 wire n_2326_o_0;
 wire n_2325_o_0;
 wire n_2324_o_0;
 wire n_2323_o_0;
 wire n_2322_o_0;
 wire n_2321_o_0;
 wire n_2320_o_0;
 wire n_2319_o_0;
 wire n_2318_o_0;
 wire n_2317_o_0;
 wire n_2316_o_0;
 wire n_2315_o_0;
 wire n_2314_o_0;
 wire n_2313_o_0;
 wire n_2312_o_0;
 wire n_2311_o_0;
 wire n_2310_o_0;
 wire n_2309_o_0;
 wire n_2308_o_0;
 wire n_2307_o_0;
 wire n_2306_o_0;
 wire n_2305_o_0;
 wire n_2304_o_0;
 wire n_2303_o_0;
 wire n_2302_o_0;
 wire n_2301_o_0;
 wire n_2300_o_0;
 wire n_2299_o_0;
 wire n_2298_o_0;
 wire n_2297_o_0;
 wire n_2296_o_0;
 wire n_2295_o_0;
 wire n_2294_o_0;
 wire n_2293_o_0;
 wire n_2292_o_0;
 wire n_2291_o_0;
 wire n_2290_o_0;
 wire n_2289_o_0;
 wire n_2288_o_0;
 wire n_2287_o_0;
 wire n_2286_o_0;
 wire n_2285_o_0;
 wire n_2284_o_0;
 wire n_2283_o_0;
 wire n_2282_o_0;
 wire n_2281_o_0;
 wire n_2280_o_0;
 wire n_2279_o_0;
 wire n_2278_o_0;
 wire n_2277_o_0;
 wire n_2276_o_0;
 wire n_2275_o_0;
 wire n_2274_o_0;
 wire n_2273_o_0;
 wire n_2272_o_0;
 wire n_2271_o_0;
 wire n_2270_o_0;
 wire n_2269_o_0;
 wire n_2268_o_0;
 wire n_2267_o_0;
 wire n_2266_o_0;
 wire n_2265_o_0;
 wire n_2264_o_0;
 wire n_2263_o_0;
 wire n_2262_o_0;
 wire n_2261_o_0;
 wire n_2260_o_0;
 wire n_2259_o_0;
 wire n_2258_o_0;
 wire n_2257_o_0;
 wire n_2256_o_0;
 wire n_2255_o_0;
 wire n_2254_o_0;
 wire n_2253_o_0;
 wire n_2252_o_0;
 wire n_2251_o_0;
 wire n_2250_o_0;
 wire n_2249_o_0;
 wire n_2248_o_0;
 wire n_2247_o_0;
 wire n_2246_o_0;
 wire n_2245_o_0;
 wire n_2244_o_0;
 wire n_2243_o_0;
 wire n_2242_o_0;
 wire n_2241_o_0;
 wire n_2240_o_0;
 wire n_2239_o_0;
 wire n_2238_o_0;
 wire n_2237_o_0;
 wire n_2236_o_0;
 wire n_2235_o_0;
 wire n_2234_o_0;
 wire n_2233_o_0;
 wire n_2232_o_0;
 wire n_2231_o_0;
 wire n_2230_o_0;
 wire n_2229_o_0;
 wire n_2228_o_0;
 wire n_2227_o_0;
 wire n_2226_o_0;
 wire n_2225_o_0;
 wire n_2224_o_0;
 wire n_2223_o_0;
 wire n_2222_o_0;
 wire n_2221_o_0;
 wire n_2220_o_0;
 wire n_2219_o_0;
 wire n_2218_o_0;
 wire n_2217_o_0;
 wire n_2216_o_0;
 wire n_2215_o_0;
 wire n_2214_o_0;
 wire n_2213_o_0;
 wire n_2212_o_0;
 wire n_2211_o_0;
 wire n_2210_o_0;
 wire n_2209_o_0;
 wire n_2208_o_0;
 wire n_2207_o_0;
 wire n_2206_o_0;
 wire n_2205_o_0;
 wire n_2204_o_0;
 wire n_2203_o_0;
 wire n_2202_o_0;
 wire n_2201_o_0;
 wire n_2200_o_0;
 wire n_2199_o_0;
 wire n_2198_o_0;
 wire n_2197_o_0;
 wire n_2196_o_0;
 wire n_2195_o_0;
 wire n_2194_o_0;
 wire n_2193_o_0;
 wire n_2192_o_0;
 wire n_2191_o_0;
 wire n_2190_o_0;
 wire n_2189_o_0;
 wire n_2188_o_0;
 wire n_2187_o_0;
 wire n_2186_o_0;
 wire n_2185_o_0;
 wire n_2184_o_0;
 wire n_2183_o_0;
 wire n_2182_o_0;
 wire n_2181_o_0;
 wire n_2180_o_0;
 wire n_2179_o_0;
 wire n_2178_o_0;
 wire n_2177_o_0;
 wire n_2176_o_0;
 wire n_2175_o_0;
 wire n_2174_o_0;
 wire n_2173_o_0;
 wire n_2172_o_0;
 wire n_2171_o_0;
 wire n_2170_o_0;
 wire n_2169_o_0;
 wire n_2168_o_0;
 wire n_2167_o_0;
 wire n_2166_o_0;
 wire n_2165_o_0;
 wire n_2164_o_0;
 wire n_2163_o_0;
 wire n_2162_o_0;
 wire n_2161_o_0;
 wire n_2160_o_0;
 wire n_2159_o_0;
 wire n_2158_o_0;
 wire n_2157_o_0;
 wire n_2156_o_0;
 wire n_2155_o_0;
 wire n_2154_o_0;
 wire n_2153_o_0;
 wire n_2152_o_0;
 wire n_2151_o_0;
 wire n_2150_o_0;
 wire n_2149_o_0;
 wire n_2148_o_0;
 wire n_2147_o_0;
 wire n_2146_o_0;
 wire n_2145_o_0;
 wire n_2144_o_0;
 wire n_2143_o_0;
 wire n_2142_o_0;
 wire n_2141_o_0;
 wire n_2140_o_0;
 wire n_2139_o_0;
 wire n_2138_o_0;
 wire n_2137_o_0;
 wire n_2136_o_0;
 wire n_2135_o_0;
 wire n_2134_o_0;
 wire n_2133_o_0;
 wire n_2132_o_0;
 wire n_2131_o_0;
 wire n_2130_o_0;
 wire n_2129_o_0;
 wire n_2128_o_0;
 wire n_2127_o_0;
 wire n_2126_o_0;
 wire n_2125_o_0;
 wire n_2124_o_0;
 wire n_2123_o_0;
 wire n_2122_o_0;
 wire n_2121_o_0;
 wire n_2120_o_0;
 wire n_2119_o_0;
 wire n_2118_o_0;
 wire n_2117_o_0;
 wire n_2116_o_0;
 wire n_2115_o_0;
 wire n_2114_o_0;
 wire n_2113_o_0;
 wire n_2112_o_0;
 wire n_2111_o_0;
 wire n_2110_o_0;
 wire n_2109_o_0;
 wire n_2108_o_0;
 wire n_2107_o_0;
 wire n_2106_o_0;
 wire n_2105_o_0;
 wire n_2104_o_0;
 wire n_2103_o_0;
 wire n_2102_o_0;
 wire n_2101_o_0;
 wire n_2100_o_0;
 wire n_2099_o_0;
 wire n_2098_o_0;
 wire n_2097_o_0;
 wire n_2096_o_0;
 wire n_2095_o_0;
 wire n_2094_o_0;
 wire n_2093_o_0;
 wire n_2092_o_0;
 wire n_2091_o_0;
 wire n_2090_o_0;
 wire n_2089_o_0;
 wire n_2088_o_0;
 wire n_2087_o_0;
 wire n_2086_o_0;
 wire n_2085_o_0;
 wire n_2084_o_0;
 wire n_2083_o_0;
 wire n_2082_o_0;
 wire n_2081_o_0;
 wire n_2080_o_0;
 wire n_2079_o_0;
 wire n_2078_o_0;
 wire n_2077_o_0;
 wire n_2076_o_0;
 wire n_2075_o_0;
 wire n_2074_o_0;
 wire n_2073_o_0;
 wire n_2072_o_0;
 wire n_2071_o_0;
 wire n_2070_o_0;
 wire n_2069_o_0;
 wire n_2068_o_0;
 wire n_2067_o_0;
 wire n_2066_o_0;
 wire n_2065_o_0;
 wire n_2064_o_0;
 wire n_2063_o_0;
 wire n_2062_o_0;
 wire n_2061_o_0;
 wire n_2060_o_0;
 wire n_2059_o_0;
 wire n_2058_o_0;
 wire n_2057_o_0;
 wire n_2056_o_0;
 wire n_2055_o_0;
 wire n_2054_o_0;
 wire n_2053_o_0;
 wire n_2052_o_0;
 wire n_2051_o_0;
 wire n_2050_o_0;
 wire n_2049_o_0;
 wire n_2048_o_0;
 wire n_2047_o_0;
 wire n_2046_o_0;
 wire n_2045_o_0;
 wire n_2044_o_0;
 wire n_2043_o_0;
 wire n_2042_o_0;
 wire n_2041_o_0;
 wire n_2040_o_0;
 wire n_2039_o_0;
 wire n_2038_o_0;
 wire n_2037_o_0;
 wire n_2036_o_0;
 wire n_2035_o_0;
 wire n_2034_o_0;
 wire n_2033_o_0;
 wire n_2032_o_0;
 wire n_2031_o_0;
 wire n_2030_o_0;
 wire n_2029_o_0;
 wire n_2028_o_0;
 wire n_2027_o_0;
 wire n_2026_o_0;
 wire n_2025_o_0;
 wire n_2024_o_0;
 wire n_2023_o_0;
 wire n_2022_o_0;
 wire n_2021_o_0;
 wire n_2020_o_0;
 wire n_2019_o_0;
 wire n_2018_o_0;
 wire n_2017_o_0;
 wire n_2016_o_0;
 wire n_2015_o_0;
 wire n_2014_o_0;
 wire n_2013_o_0;
 wire n_2012_o_0;
 wire n_2011_o_0;
 wire n_2010_o_0;
 wire n_2009_o_0;
 wire n_2008_o_0;
 wire n_2007_o_0;
 wire n_2006_o_0;
 wire n_2005_o_0;
 wire n_2004_o_0;
 wire n_2003_o_0;
 wire n_2002_o_0;
 wire n_2001_o_0;
 wire n_2000_o_0;
 wire n_1999_o_0;
 wire n_1998_o_0;
 wire n_1997_o_0;
 wire n_1996_o_0;
 wire n_1995_o_0;
 wire n_1994_o_0;
 wire n_1993_o_0;
 wire n_1992_o_0;
 wire n_1991_o_0;
 wire n_1990_o_0;
 wire n_1989_o_0;
 wire n_1988_o_0;
 wire n_1987_o_0;
 wire n_1986_o_0;
 wire n_1985_o_0;
 wire n_1984_o_0;
 wire n_1983_o_0;
 wire n_1982_o_0;
 wire n_1981_o_0;
 wire n_1980_o_0;
 wire n_1979_o_0;
 wire n_1978_o_0;
 wire n_1977_o_0;
 wire n_1976_o_0;
 wire n_1975_o_0;
 wire n_1974_o_0;
 wire n_1973_o_0;
 wire n_1972_o_0;
 wire n_1971_o_0;
 wire n_1970_o_0;
 wire n_1969_o_0;
 wire n_1968_o_0;
 wire n_1967_o_0;
 wire n_1966_o_0;
 wire n_1965_o_0;
 wire n_1964_o_0;
 wire n_1963_o_0;
 wire n_1962_o_0;
 wire n_1961_o_0;
 wire n_1960_o_0;
 wire n_1959_o_0;
 wire n_1958_o_0;
 wire n_1957_o_0;
 wire n_1956_o_0;
 wire n_1955_o_0;
 wire n_1954_o_0;
 wire n_1953_o_0;
 wire n_1952_o_0;
 wire n_1951_o_0;
 wire n_1950_o_0;
 wire n_1949_o_0;
 wire n_1948_o_0;
 wire n_1947_o_0;
 wire n_1946_o_0;
 wire n_1945_o_0;
 wire n_1944_o_0;
 wire n_1943_o_0;
 wire n_1942_o_0;
 wire n_1941_o_0;
 wire n_1940_o_0;
 wire n_1939_o_0;
 wire n_1938_o_0;
 wire n_1937_o_0;
 wire n_1936_o_0;
 wire n_1935_o_0;
 wire n_1934_o_0;
 wire n_1933_o_0;
 wire n_1932_o_0;
 wire n_1931_o_0;
 wire n_1930_o_0;
 wire n_1929_o_0;
 wire n_1928_o_0;
 wire n_1927_o_0;
 wire n_1926_o_0;
 wire n_1925_o_0;
 wire n_1924_o_0;
 wire n_1923_o_0;
 wire n_1922_o_0;
 wire n_1921_o_0;
 wire n_1920_o_0;
 wire n_1919_o_0;
 wire n_1918_o_0;
 wire n_1917_o_0;
 wire n_1916_o_0;
 wire n_1915_o_0;
 wire n_1914_o_0;
 wire n_1913_o_0;
 wire n_1912_o_0;
 wire n_1911_o_0;
 wire n_1910_o_0;
 wire n_1909_o_0;
 wire n_1908_o_0;
 wire n_1907_o_0;
 wire n_1906_o_0;
 wire n_1905_o_0;
 wire n_1904_o_0;
 wire n_1903_o_0;
 wire n_1902_o_0;
 wire n_1901_o_0;
 wire n_1900_o_0;
 wire n_1899_o_0;
 wire n_1898_o_0;
 wire n_1897_o_0;
 wire n_1896_o_0;
 wire n_1895_o_0;
 wire n_1894_o_0;
 wire n_1893_o_0;
 wire n_1892_o_0;
 wire n_1891_o_0;
 wire n_1890_o_0;
 wire n_1889_o_0;
 wire n_1888_o_0;
 wire n_1887_o_0;
 wire n_1886_o_0;
 wire n_1885_o_0;
 wire n_1884_o_0;
 wire n_1883_o_0;
 wire n_1882_o_0;
 wire n_1881_o_0;
 wire n_1880_o_0;
 wire n_1879_o_0;
 wire n_1878_o_0;
 wire n_1877_o_0;
 wire n_1876_o_0;
 wire n_1875_o_0;
 wire n_1874_o_0;
 wire n_1873_o_0;
 wire n_1872_o_0;
 wire n_1871_o_0;
 wire n_1870_o_0;
 wire n_1869_o_0;
 wire n_1868_o_0;
 wire n_1867_o_0;
 wire n_1866_o_0;
 wire n_1865_o_0;
 wire n_1864_o_0;
 wire n_1863_o_0;
 wire n_1862_o_0;
 wire n_1861_o_0;
 wire n_1860_o_0;
 wire n_1859_o_0;
 wire n_1858_o_0;
 wire n_1857_o_0;
 wire n_1856_o_0;
 wire n_1855_o_0;
 wire n_1854_o_0;
 wire n_1853_o_0;
 wire n_1852_o_0;
 wire n_1851_o_0;
 wire n_1850_o_0;
 wire n_1849_o_0;
 wire n_1848_o_0;
 wire n_1847_o_0;
 wire n_1846_o_0;
 wire n_1845_o_0;
 wire n_1844_o_0;
 wire n_1843_o_0;
 wire n_1842_o_0;
 wire n_1841_o_0;
 wire n_1840_o_0;
 wire n_1839_o_0;
 wire n_1838_o_0;
 wire n_1837_o_0;
 wire n_1836_o_0;
 wire n_1835_o_0;
 wire n_1834_o_0;
 wire n_1833_o_0;
 wire n_1832_o_0;
 wire n_1831_o_0;
 wire n_1830_o_0;
 wire n_1829_o_0;
 wire n_1828_o_0;
 wire n_1827_o_0;
 wire n_1826_o_0;
 wire n_1825_o_0;
 wire n_1824_o_0;
 wire n_1823_o_0;
 wire n_1822_o_0;
 wire n_1821_o_0;
 wire n_1820_o_0;
 wire n_1819_o_0;
 wire n_1818_o_0;
 wire n_1817_o_0;
 wire n_1816_o_0;
 wire n_1815_o_0;
 wire n_1814_o_0;
 wire n_1813_o_0;
 wire n_1812_o_0;
 wire n_1811_o_0;
 wire n_1810_o_0;
 wire n_1809_o_0;
 wire n_1808_o_0;
 wire n_1807_o_0;
 wire n_1806_o_0;
 wire n_1805_o_0;
 wire n_1804_o_0;
 wire n_1803_o_0;
 wire n_1802_o_0;
 wire n_1801_o_0;
 wire n_1800_o_0;
 wire n_1799_o_0;
 wire n_1798_o_0;
 wire n_1797_o_0;
 wire n_1796_o_0;
 wire n_1795_o_0;
 wire n_1794_o_0;
 wire n_1793_o_0;
 wire n_1792_o_0;
 wire n_1791_o_0;
 wire n_1790_o_0;
 wire n_1789_o_0;
 wire n_1788_o_0;
 wire n_1787_o_0;
 wire n_1786_o_0;
 wire n_1785_o_0;
 wire n_1784_o_0;
 wire n_1783_o_0;
 wire n_1782_o_0;
 wire n_1781_o_0;
 wire n_1780_o_0;
 wire n_1779_o_0;
 wire n_1778_o_0;
 wire n_1777_o_0;
 wire n_1776_o_0;
 wire n_1775_o_0;
 wire n_1774_o_0;
 wire n_1773_o_0;
 wire n_1772_o_0;
 wire n_1771_o_0;
 wire n_1770_o_0;
 wire n_1769_o_0;
 wire n_1768_o_0;
 wire n_1767_o_0;
 wire n_1766_o_0;
 wire n_1765_o_0;
 wire n_1764_o_0;
 wire n_1763_o_0;
 wire n_1762_o_0;
 wire n_1761_o_0;
 wire n_1760_o_0;
 wire n_1759_o_0;
 wire n_1758_o_0;
 wire n_1757_o_0;
 wire n_1756_o_0;
 wire n_1755_o_0;
 wire n_1754_o_0;
 wire n_1753_o_0;
 wire n_1752_o_0;
 wire n_1751_o_0;
 wire n_1750_o_0;
 wire n_1749_o_0;
 wire n_1748_o_0;
 wire n_1747_o_0;
 wire n_1746_o_0;
 wire n_1745_o_0;
 wire n_1744_o_0;
 wire n_1743_o_0;
 wire n_1742_o_0;
 wire n_1741_o_0;
 wire n_1740_o_0;
 wire n_1739_o_0;
 wire n_1738_o_0;
 wire n_1737_o_0;
 wire n_1736_o_0;
 wire n_1735_o_0;
 wire n_1734_o_0;
 wire n_1733_o_0;
 wire n_1732_o_0;
 wire n_1731_o_0;
 wire n_1730_o_0;
 wire n_1729_o_0;
 wire n_1728_o_0;
 wire n_1727_o_0;
 wire n_1726_o_0;
 wire n_1725_o_0;
 wire n_1724_o_0;
 wire n_1723_o_0;
 wire n_1722_o_0;
 wire n_1721_o_0;
 wire n_1720_o_0;
 wire n_1719_o_0;
 wire n_1718_o_0;
 wire n_1717_o_0;
 wire n_1716_o_0;
 wire n_1715_o_0;
 wire n_1714_o_0;
 wire n_1713_o_0;
 wire n_1712_o_0;
 wire n_1711_o_0;
 wire n_1710_o_0;
 wire n_1709_o_0;
 wire n_1708_o_0;
 wire n_1707_o_0;
 wire n_1706_o_0;
 wire n_1705_o_0;
 wire n_1704_o_0;
 wire n_1703_o_0;
 wire n_1702_o_0;
 wire n_1701_o_0;
 wire n_1700_o_0;
 wire n_1699_o_0;
 wire n_1698_o_0;
 wire n_1697_o_0;
 wire n_1696_o_0;
 wire n_1695_o_0;
 wire n_1694_o_0;
 wire n_1693_o_0;
 wire n_1692_o_0;
 wire n_1691_o_0;
 wire n_1690_o_0;
 wire n_1689_o_0;
 wire n_1688_o_0;
 wire n_1687_o_0;
 wire n_1686_o_0;
 wire n_1685_o_0;
 wire n_1684_o_0;
 wire n_1683_o_0;
 wire n_1682_o_0;
 wire n_1681_o_0;
 wire n_1680_o_0;
 wire n_1679_o_0;
 wire n_1678_o_0;
 wire n_1677_o_0;
 wire n_1676_o_0;
 wire n_1675_o_0;
 wire n_1674_o_0;
 wire n_1673_o_0;
 wire n_1672_o_0;
 wire n_1671_o_0;
 wire n_1670_o_0;
 wire n_1669_o_0;
 wire n_1668_o_0;
 wire n_1667_o_0;
 wire n_1666_o_0;
 wire n_1665_o_0;
 wire n_1664_o_0;
 wire n_1663_o_0;
 wire n_1662_o_0;
 wire n_1661_o_0;
 wire n_1660_o_0;
 wire n_1659_o_0;
 wire n_1658_o_0;
 wire n_1657_o_0;
 wire n_1656_o_0;
 wire n_1655_o_0;
 wire n_1654_o_0;
 wire n_1653_o_0;
 wire n_1652_o_0;
 wire n_1651_o_0;
 wire n_1650_o_0;
 wire n_1649_o_0;
 wire n_1648_o_0;
 wire n_1647_o_0;
 wire n_1646_o_0;
 wire n_1645_o_0;
 wire n_1644_o_0;
 wire n_1643_o_0;
 wire n_1642_o_0;
 wire n_1641_o_0;
 wire n_1640_o_0;
 wire n_1639_o_0;
 wire n_1638_o_0;
 wire n_1637_o_0;
 wire n_1636_o_0;
 wire n_1635_o_0;
 wire n_1634_o_0;
 wire n_1633_o_0;
 wire n_1632_o_0;
 wire n_1631_o_0;
 wire n_1630_o_0;
 wire n_1629_o_0;
 wire n_1628_o_0;
 wire n_1627_o_0;
 wire n_1626_o_0;
 wire n_1625_o_0;
 wire n_1624_o_0;
 wire n_1623_o_0;
 wire n_1622_o_0;
 wire n_1621_o_0;
 wire n_1620_o_0;
 wire n_1619_o_0;
 wire n_1618_o_0;
 wire n_1617_o_0;
 wire n_1616_o_0;
 wire n_1615_o_0;
 wire n_1614_o_0;
 wire n_1613_o_0;
 wire n_1612_o_0;
 wire n_1611_o_0;
 wire n_1610_o_0;
 wire n_1609_o_0;
 wire n_1608_o_0;
 wire n_1607_o_0;
 wire n_1606_o_0;
 wire n_1605_o_0;
 wire n_1604_o_0;
 wire n_1603_o_0;
 wire n_1602_o_0;
 wire n_1601_o_0;
 wire n_1600_o_0;
 wire n_1599_o_0;
 wire n_1598_o_0;
 wire n_1597_o_0;
 wire n_1596_o_0;
 wire n_1595_o_0;
 wire n_1594_o_0;
 wire n_1593_o_0;
 wire n_1592_o_0;
 wire n_1591_o_0;
 wire n_1590_o_0;
 wire n_1589_o_0;
 wire n_1588_o_0;
 wire n_1587_o_0;
 wire n_1586_o_0;
 wire n_1585_o_0;
 wire n_1584_o_0;
 wire n_1583_o_0;
 wire n_1582_o_0;
 wire n_1581_o_0;
 wire n_1580_o_0;
 wire n_1579_o_0;
 wire n_1578_o_0;
 wire n_1577_o_0;
 wire n_1576_o_0;
 wire n_1575_o_0;
 wire n_1574_o_0;
 wire n_1573_o_0;
 wire n_1572_o_0;
 wire n_1571_o_0;
 wire n_1570_o_0;
 wire n_1569_o_0;
 wire n_1568_o_0;
 wire n_1567_o_0;
 wire n_1566_o_0;
 wire n_1565_o_0;
 wire n_1564_o_0;
 wire n_1563_o_0;
 wire n_1562_o_0;
 wire n_1561_o_0;
 wire n_1560_o_0;
 wire n_1559_o_0;
 wire n_1558_o_0;
 wire n_1557_o_0;
 wire n_1556_o_0;
 wire n_1555_o_0;
 wire n_1554_o_0;
 wire n_1553_o_0;
 wire n_1552_o_0;
 wire n_1551_o_0;
 wire n_1550_o_0;
 wire n_1549_o_0;
 wire n_1548_o_0;
 wire n_1547_o_0;
 wire n_1546_o_0;
 wire n_1545_o_0;
 wire n_1544_o_0;
 wire n_1543_o_0;
 wire n_1542_o_0;
 wire n_1541_o_0;
 wire n_1540_o_0;
 wire n_1539_o_0;
 wire n_1538_o_0;
 wire n_1537_o_0;
 wire n_1536_o_0;
 wire n_1535_o_0;
 wire n_1534_o_0;
 wire n_1533_o_0;
 wire n_1532_o_0;
 wire n_1531_o_0;
 wire n_1530_o_0;
 wire n_1529_o_0;
 wire n_1528_o_0;
 wire n_1527_o_0;
 wire n_1526_o_0;
 wire n_1525_o_0;
 wire n_1524_o_0;
 wire n_1523_o_0;
 wire n_1522_o_0;
 wire n_1521_o_0;
 wire n_1520_o_0;
 wire n_1519_o_0;
 wire n_1518_o_0;
 wire n_1517_o_0;
 wire n_1516_o_0;
 wire n_1515_o_0;
 wire n_1514_o_0;
 wire n_1513_o_0;
 wire n_1512_o_0;
 wire n_1511_o_0;
 wire n_1510_o_0;
 wire n_1509_o_0;
 wire n_1508_o_0;
 wire n_1507_o_0;
 wire n_1506_o_0;
 wire n_1505_o_0;
 wire n_1504_o_0;
 wire n_1503_o_0;
 wire n_1502_o_0;
 wire n_1501_o_0;
 wire n_1500_o_0;
 wire n_1499_o_0;
 wire n_1498_o_0;
 wire n_1497_o_0;
 wire n_1496_o_0;
 wire n_1495_o_0;
 wire n_1494_o_0;
 wire n_1493_o_0;
 wire n_1492_o_0;
 wire n_1491_o_0;
 wire n_1490_o_0;
 wire n_1489_o_0;
 wire n_1488_o_0;
 wire n_1487_o_0;
 wire n_1486_o_0;
 wire n_1485_o_0;
 wire n_1484_o_0;
 wire n_1483_o_0;
 wire n_1482_o_0;
 wire n_1481_o_0;
 wire n_1480_o_0;
 wire n_1479_o_0;
 wire n_1478_o_0;
 wire n_1477_o_0;
 wire n_1476_o_0;
 wire n_1475_o_0;
 wire n_1474_o_0;
 wire n_1473_o_0;
 wire n_1472_o_0;
 wire n_1471_o_0;
 wire n_1470_o_0;
 wire n_1469_o_0;
 wire n_1468_o_0;
 wire n_1467_o_0;
 wire n_1466_o_0;
 wire n_1465_o_0;
 wire n_1464_o_0;
 wire n_1463_o_0;
 wire n_1462_o_0;
 wire n_1461_o_0;
 wire n_1460_o_0;
 wire n_1459_o_0;
 wire n_1458_o_0;
 wire n_1457_o_0;
 wire n_1456_o_0;
 wire n_1455_o_0;
 wire n_1454_o_0;
 wire n_1453_o_0;
 wire n_1452_o_0;
 wire n_1451_o_0;
 wire n_1450_o_0;
 wire n_1449_o_0;
 wire n_1448_o_0;
 wire n_1447_o_0;
 wire n_1446_o_0;
 wire n_1445_o_0;
 wire n_1444_o_0;
 wire n_1443_o_0;
 wire n_1442_o_0;
 wire n_1441_o_0;
 wire n_1440_o_0;
 wire n_1439_o_0;
 wire n_1438_o_0;
 wire n_1437_o_0;
 wire n_1436_o_0;
 wire n_1435_o_0;
 wire n_1434_o_0;
 wire n_1433_o_0;
 wire n_1432_o_0;
 wire n_1431_o_0;
 wire n_1430_o_0;
 wire n_1429_o_0;
 wire n_1428_o_0;
 wire n_1427_o_0;
 wire n_1426_o_0;
 wire n_1425_o_0;
 wire n_1424_o_0;
 wire n_1423_o_0;
 wire n_1422_o_0;
 wire n_1421_o_0;
 wire n_1420_o_0;
 wire n_1419_o_0;
 wire n_1418_o_0;
 wire n_1417_o_0;
 wire n_1416_o_0;
 wire n_1415_o_0;
 wire n_1414_o_0;
 wire n_1413_o_0;
 wire n_1412_o_0;
 wire n_1411_o_0;
 wire n_1410_o_0;
 wire n_1409_o_0;
 wire n_1408_o_0;
 wire n_1407_o_0;
 wire n_1406_o_0;
 wire n_1405_o_0;
 wire n_1404_o_0;
 wire n_1403_o_0;
 wire n_1402_o_0;
 wire n_1401_o_0;
 wire n_1400_o_0;
 wire n_1399_o_0;
 wire n_1398_o_0;
 wire n_1397_o_0;
 wire n_1396_o_0;
 wire n_1395_o_0;
 wire n_1394_o_0;
 wire n_1393_o_0;
 wire n_1392_o_0;
 wire n_1391_o_0;
 wire n_1390_o_0;
 wire n_1389_o_0;
 wire n_1388_o_0;
 wire n_1387_o_0;
 wire n_1386_o_0;
 wire n_1385_o_0;
 wire n_1384_o_0;
 wire n_1383_o_0;
 wire n_1382_o_0;
 wire n_1381_o_0;
 wire n_1380_o_0;
 wire n_1379_o_0;
 wire n_1378_o_0;
 wire n_1377_o_0;
 wire n_1376_o_0;
 wire n_1375_o_0;
 wire n_1374_o_0;
 wire n_1373_o_0;
 wire n_1372_o_0;
 wire n_1371_o_0;
 wire n_1370_o_0;
 wire n_1369_o_0;
 wire n_1368_o_0;
 wire n_1367_o_0;
 wire n_1366_o_0;
 wire n_1365_o_0;
 wire n_1364_o_0;
 wire n_1363_o_0;
 wire n_1362_o_0;
 wire n_1361_o_0;
 wire n_1360_o_0;
 wire n_1359_o_0;
 wire n_1358_o_0;
 wire n_1357_o_0;
 wire n_1356_o_0;
 wire n_1355_o_0;
 wire n_1354_o_0;
 wire n_1353_o_0;
 wire n_1352_o_0;
 wire n_1351_o_0;
 wire n_1350_o_0;
 wire n_1349_o_0;
 wire n_1348_o_0;
 wire n_1347_o_0;
 wire n_1346_o_0;
 wire n_1345_o_0;
 wire n_1344_o_0;
 wire n_1343_o_0;
 wire n_1342_o_0;
 wire n_1341_o_0;
 wire n_1340_o_0;
 wire n_1339_o_0;
 wire n_1338_o_0;
 wire n_1337_o_0;
 wire n_1336_o_0;
 wire n_1335_o_0;
 wire n_1334_o_0;
 wire n_1333_o_0;
 wire n_1332_o_0;
 wire n_1331_o_0;
 wire n_1330_o_0;
 wire n_1329_o_0;
 wire n_1328_o_0;
 wire n_1327_o_0;
 wire n_1326_o_0;
 wire n_1325_o_0;
 wire n_1324_o_0;
 wire n_1323_o_0;
 wire n_1322_o_0;
 wire n_1321_o_0;
 wire n_1320_o_0;
 wire n_1319_o_0;
 wire n_1318_o_0;
 wire n_1317_o_0;
 wire n_1316_o_0;
 wire n_1315_o_0;
 wire n_1314_o_0;
 wire n_1313_o_0;
 wire n_1312_o_0;
 wire n_1311_o_0;
 wire n_1310_o_0;
 wire n_1309_o_0;
 wire n_1308_o_0;
 wire n_1307_o_0;
 wire n_1306_o_0;
 wire n_1305_o_0;
 wire n_1304_o_0;
 wire n_1303_o_0;
 wire n_1302_o_0;
 wire n_1301_o_0;
 wire n_1300_o_0;
 wire n_1299_o_0;
 wire n_1298_o_0;
 wire n_1297_o_0;
 wire n_1296_o_0;
 wire n_1295_o_0;
 wire n_1294_o_0;
 wire n_1293_o_0;
 wire n_1292_o_0;
 wire n_1291_o_0;
 wire n_1290_o_0;
 wire n_1289_o_0;
 wire n_1288_o_0;
 wire n_1287_o_0;
 wire n_1286_o_0;
 wire n_1285_o_0;
 wire n_1284_o_0;
 wire n_1283_o_0;
 wire n_1282_o_0;
 wire n_1281_o_0;
 wire n_1280_o_0;
 wire n_1279_o_0;
 wire n_1278_o_0;
 wire n_1277_o_0;
 wire n_1276_o_0;
 wire n_1275_o_0;
 wire n_1274_o_0;
 wire n_1273_o_0;
 wire n_1272_o_0;
 wire n_1271_o_0;
 wire n_1270_o_0;
 wire n_1269_o_0;
 wire n_1268_o_0;
 wire n_1267_o_0;
 wire n_1266_o_0;
 wire n_1265_o_0;
 wire n_1264_o_0;
 wire n_1263_o_0;
 wire n_1262_o_0;
 wire n_1261_o_0;
 wire n_1260_o_0;
 wire n_1259_o_0;
 wire n_1258_o_0;
 wire n_1257_o_0;
 wire n_1256_o_0;
 wire n_1255_o_0;
 wire n_1254_o_0;
 wire n_1253_o_0;
 wire n_1252_o_0;
 wire n_1251_o_0;
 wire n_1250_o_0;
 wire n_1249_o_0;
 wire n_1248_o_0;
 wire n_1247_o_0;
 wire n_1246_o_0;
 wire n_1245_o_0;
 wire n_1244_o_0;
 wire n_1243_o_0;
 wire n_1242_o_0;
 wire n_1241_o_0;
 wire n_1240_o_0;
 wire n_1239_o_0;
 wire n_1238_o_0;
 wire n_1237_o_0;
 wire n_1236_o_0;
 wire n_1235_o_0;
 wire n_1234_o_0;
 wire n_1233_o_0;
 wire n_1232_o_0;
 wire n_1231_o_0;
 wire n_1230_o_0;
 wire n_1229_o_0;
 wire n_1228_o_0;
 wire n_1227_o_0;
 wire n_1226_o_0;
 wire n_1225_o_0;
 wire n_1224_o_0;
 wire n_1223_o_0;
 wire n_1222_o_0;
 wire n_1221_o_0;
 wire n_1220_o_0;
 wire n_1219_o_0;
 wire n_1218_o_0;
 wire n_1217_o_0;
 wire n_1216_o_0;
 wire n_1215_o_0;
 wire n_1214_o_0;
 wire n_1213_o_0;
 wire n_1212_o_0;
 wire n_1211_o_0;
 wire n_1210_o_0;
 wire n_1209_o_0;
 wire n_1208_o_0;
 wire n_1207_o_0;
 wire n_1206_o_0;
 wire n_1205_o_0;
 wire n_1204_o_0;
 wire n_1203_o_0;
 wire n_1202_o_0;
 wire n_1201_o_0;
 wire n_1200_o_0;
 wire n_1199_o_0;
 wire n_1198_o_0;
 wire n_1197_o_0;
 wire n_1196_o_0;
 wire n_1195_o_0;
 wire n_1194_o_0;
 wire n_1193_o_0;
 wire n_1192_o_0;
 wire n_1191_o_0;
 wire n_1190_o_0;
 wire n_1189_o_0;
 wire n_1188_o_0;
 wire n_1187_o_0;
 wire n_1186_o_0;
 wire n_1185_o_0;
 wire n_1184_o_0;
 wire n_1183_o_0;
 wire n_1182_o_0;
 wire n_1181_o_0;
 wire n_1180_o_0;
 wire n_1179_o_0;
 wire n_1178_o_0;
 wire n_1177_o_0;
 wire n_1176_o_0;
 wire n_1175_o_0;
 wire n_1174_o_0;
 wire n_1173_o_0;
 wire n_1172_o_0;
 wire n_1171_o_0;
 wire n_1170_o_0;
 wire n_1169_o_0;
 wire n_1168_o_0;
 wire n_1167_o_0;
 wire n_1166_o_0;
 wire n_1165_o_0;
 wire n_1164_o_0;
 wire n_1163_o_0;
 wire n_1162_o_0;
 wire n_1161_o_0;
 wire n_1160_o_0;
 wire n_1159_o_0;
 wire n_1158_o_0;
 wire n_1157_o_0;
 wire n_1156_o_0;
 wire n_1155_o_0;
 wire n_1154_o_0;
 wire n_1153_o_0;
 wire n_1152_o_0;
 wire n_1151_o_0;
 wire n_1150_o_0;
 wire n_1149_o_0;
 wire n_1148_o_0;
 wire n_1147_o_0;
 wire n_1146_o_0;
 wire n_1145_o_0;
 wire n_1144_o_0;
 wire n_1143_o_0;
 wire n_1142_o_0;
 wire n_1141_o_0;
 wire n_1140_o_0;
 wire n_1139_o_0;
 wire n_1138_o_0;
 wire n_1137_o_0;
 wire n_1136_o_0;
 wire n_1135_o_0;
 wire n_1134_o_0;
 wire n_1133_o_0;
 wire n_1132_o_0;
 wire n_1131_o_0;
 wire n_1130_o_0;
 wire n_1129_o_0;
 wire n_1128_o_0;
 wire n_1127_o_0;
 wire n_1126_o_0;
 wire n_1125_o_0;
 wire n_1124_o_0;
 wire n_1123_o_0;
 wire n_1122_o_0;
 wire n_1121_o_0;
 wire n_1120_o_0;
 wire n_1119_o_0;
 wire n_1118_o_0;
 wire n_1117_o_0;
 wire n_1116_o_0;
 wire n_1115_o_0;
 wire n_1114_o_0;
 wire n_1113_o_0;
 wire n_1112_o_0;
 wire n_1111_o_0;
 wire n_1110_o_0;
 wire n_1109_o_0;
 wire n_1108_o_0;
 wire n_1107_o_0;
 wire n_1106_o_0;
 wire n_1105_o_0;
 wire n_1104_o_0;
 wire n_1103_o_0;
 wire n_1102_o_0;
 wire n_1101_o_0;
 wire n_1100_o_0;
 wire n_1099_o_0;
 wire n_1098_o_0;
 wire n_1097_o_0;
 wire n_1096_o_0;
 wire n_1095_o_0;
 wire n_1094_o_0;
 wire n_1093_o_0;
 wire n_1092_o_0;
 wire n_1091_o_0;
 wire n_1090_o_0;
 wire n_1089_o_0;
 wire n_1088_o_0;
 wire n_1087_o_0;
 wire n_1086_o_0;
 wire n_1085_o_0;
 wire n_1084_o_0;
 wire n_1083_o_0;
 wire n_1082_o_0;
 wire n_1081_o_0;
 wire n_1080_o_0;
 wire n_1079_o_0;
 wire n_1078_o_0;
 wire n_1077_o_0;
 wire n_1076_o_0;
 wire n_1075_o_0;
 wire n_1074_o_0;
 wire n_1073_o_0;
 wire n_1072_o_0;
 wire n_1071_o_0;
 wire n_1070_o_0;
 wire n_1069_o_0;
 wire n_1068_o_0;
 wire n_1067_o_0;
 wire n_1066_o_0;
 wire n_1065_o_0;
 wire n_1064_o_0;
 wire n_1063_o_0;
 wire n_1062_o_0;
 wire n_1061_o_0;
 wire n_1060_o_0;
 wire n_1059_o_0;
 wire n_1058_o_0;
 wire n_1057_o_0;
 wire n_1056_o_0;
 wire n_1055_o_0;
 wire n_1054_o_0;
 wire n_1053_o_0;
 wire n_1052_o_0;
 wire n_1051_o_0;
 wire n_1050_o_0;
 wire n_1049_o_0;
 wire n_1048_o_0;
 wire n_1047_o_0;
 wire n_1046_o_0;
 wire n_1045_o_0;
 wire n_1044_o_0;
 wire n_1043_o_0;
 wire n_1042_o_0;
 wire n_1041_o_0;
 wire n_1040_o_0;
 wire n_1039_o_0;
 wire n_1038_o_0;
 wire n_1037_o_0;
 wire n_1036_o_0;
 wire n_1035_o_0;
 wire n_1034_o_0;
 wire n_1033_o_0;
 wire n_1032_o_0;
 wire n_1031_o_0;
 wire n_1030_o_0;
 wire n_1029_o_0;
 wire n_1028_o_0;
 wire n_1027_o_0;
 wire n_1026_o_0;
 wire n_1025_o_0;
 wire n_1024_o_0;
 wire n_1023_o_0;
 wire n_1022_o_0;
 wire n_1021_o_0;
 wire n_1020_o_0;
 wire n_1019_o_0;
 wire n_1018_o_0;
 wire n_1017_o_0;
 wire n_1016_o_0;
 wire n_1015_o_0;
 wire n_1014_o_0;
 wire n_1013_o_0;
 wire n_1012_o_0;
 wire n_1011_o_0;
 wire n_1010_o_0;
 wire n_1009_o_0;
 wire n_1008_o_0;
 wire n_1007_o_0;
 wire n_1006_o_0;
 wire n_1005_o_0;
 wire n_1004_o_0;
 wire n_1003_o_0;
 wire n_1002_o_0;
 wire n_1001_o_0;
 wire n_1000_o_0;
 wire n_999_o_0;
 wire n_998_o_0;
 wire n_997_o_0;
 wire n_996_o_0;
 wire n_995_o_0;
 wire n_994_o_0;
 wire n_993_o_0;
 wire n_992_o_0;
 wire n_991_o_0;
 wire n_990_o_0;
 wire n_989_o_0;
 wire n_988_o_0;
 wire n_987_o_0;
 wire n_986_o_0;
 wire n_985_o_0;
 wire n_984_o_0;
 wire n_983_o_0;
 wire n_982_o_0;
 wire n_981_o_0;
 wire n_980_o_0;
 wire n_979_o_0;
 wire n_978_o_0;
 wire n_977_o_0;
 wire n_976_o_0;
 wire n_975_o_0;
 wire n_974_o_0;
 wire n_973_o_0;
 wire n_972_o_0;
 wire n_971_o_0;
 wire n_970_o_0;
 wire n_969_o_0;
 wire n_968_o_0;
 wire n_967_o_0;
 wire n_966_o_0;
 wire n_965_o_0;
 wire n_964_o_0;
 wire n_963_o_0;
 wire n_962_o_0;
 wire n_961_o_0;
 wire n_960_o_0;
 wire n_959_o_0;
 wire n_958_o_0;
 wire n_957_o_0;
 wire n_956_o_0;
 wire n_955_o_0;
 wire n_954_o_0;
 wire n_953_o_0;
 wire n_952_o_0;
 wire n_951_o_0;
 wire n_950_o_0;
 wire n_949_o_0;
 wire n_948_o_0;
 wire n_947_o_0;
 wire n_946_o_0;
 wire n_945_o_0;
 wire n_944_o_0;
 wire n_943_o_0;
 wire n_942_o_0;
 wire n_941_o_0;
 wire n_940_o_0;
 wire n_939_o_0;
 wire n_938_o_0;
 wire n_937_o_0;
 wire n_936_o_0;
 wire n_935_o_0;
 wire n_934_o_0;
 wire n_933_o_0;
 wire n_932_o_0;
 wire n_931_o_0;
 wire _11695_;
 wire n_930_o_0;
 wire n_929_o_0;
 wire n_928_o_0;
 wire n_927_o_0;
 wire n_926_o_0;
 wire n_925_o_0;
 wire n_924_o_0;
 wire n_923_o_0;
 wire n_922_o_0;
 wire n_921_o_0;
 wire n_920_o_0;
 wire n_919_o_0;
 wire n_918_o_0;
 wire n_917_o_0;
 wire n_916_o_0;
 wire n_915_o_0;
 wire n_914_o_0;
 wire n_913_o_0;
 wire n_912_o_0;
 wire n_911_o_0;
 wire n_910_o_0;
 wire n_909_o_1;
 wire n_909_o_0;
 wire n_908_o_0;
 wire n_907_o_0;
 wire n_906_o_0;
 wire n_905_o_0;
 wire n_904_o_0;
 wire n_903_o_0;
 wire n_902_o_0;
 wire n_901_o_0;
 wire n_900_o_0;
 wire n_899_o_0;
 wire n_898_o_0;
 wire n_897_o_0;
 wire n_896_o_0;
 wire n_895_o_0;
 wire n_894_o_0;
 wire n_893_o_0;
 wire n_892_o_0;
 wire n_891_o_0;
 wire n_890_o_0;
 wire n_889_o_0;
 wire n_888_o_0;
 wire n_887_o_0;
 wire n_886_o_0;
 wire n_885_o_0;
 wire n_884_o_0;
 wire n_883_o_0;
 wire n_882_o_0;
 wire n_881_o_0;
 wire n_880_o_0;
 wire n_879_o_0;
 wire n_878_o_0;
 wire n_877_o_0;
 wire n_876_o_0;
 wire n_875_o_0;
 wire n_874_o_0;
 wire n_873_o_0;
 wire n_872_o_0;
 wire n_871_o_0;
 wire n_870_o_0;
 wire n_869_o_0;
 wire n_868_o_0;
 wire n_867_o_0;
 wire n_866_o_0;
 wire n_865_o_0;
 wire n_864_o_0;
 wire n_863_o_0;
 wire n_862_o_0;
 wire n_861_o_0;
 wire n_860_o_0;
 wire n_859_o_0;
 wire n_858_o_0;
 wire n_857_o_0;
 wire n_856_o_0;
 wire n_855_o_0;
 wire n_854_o_0;
 wire n_853_o_0;
 wire n_852_o_0;
 wire n_851_o_0;
 wire n_850_o_0;
 wire n_849_o_0;
 wire n_848_o_0;
 wire n_847_o_0;
 wire n_846_o_0;
 wire n_845_o_0;
 wire n_844_o_0;
 wire n_843_o_0;
 wire n_842_o_0;
 wire n_841_o_0;
 wire n_840_o_0;
 wire n_839_o_0;
 wire n_838_o_0;
 wire n_837_o_0;
 wire n_836_o_0;
 wire n_835_o_0;
 wire n_834_o_0;
 wire n_833_o_0;
 wire n_832_o_0;
 wire n_831_o_0;
 wire n_830_o_0;
 wire n_829_o_0;
 wire n_828_o_0;
 wire n_827_o_0;
 wire n_826_o_0;
 wire n_825_o_0;
 wire n_824_o_0;
 wire net102;
 wire net101;
 wire net100;
 wire net99;
 wire net98;
 wire net97;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net90;
 wire net89;
 wire net86;
 wire net85;
 wire net82;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire n_823_o_0;
 wire n_822_o_0;
 wire \u0/r0/rcnt_next[0] ;
 wire n_11513_o_0;
 wire n_11514_o_0;
 wire n_11515_o_0;
 wire n_11516_o_0;
 wire n_11517_o_0;
 wire n_11518_o_0;
 wire n_11519_o_0;
 wire n_11520_o_0;
 wire n_11521_o_0;
 wire n_11522_o_0;
 wire n_11523_o_0;
 wire n_11524_o_0;
 wire n_11525_o_0;
 wire n_11526_o_0;
 wire n_11527_o_0;
 wire n_11528_o_0;
 wire n_11529_o_0;
 wire n_11530_o_0;
 wire n_11531_o_0;
 wire n_11532_o_0;
 wire n_11533_o_0;
 wire n_11534_o_0;
 wire n_11535_o_0;
 wire n_11536_o_0;
 wire n_11537_o_0;
 wire n_11538_o_0;
 wire n_11539_o_0;
 wire n_11540_o_0;
 wire n_11541_o_0;
 wire n_11542_o_0;
 wire n_11543_o_0;
 wire n_11544_o_0;
 wire n_11545_o_0;
 wire n_11546_o_0;
 wire n_11547_o_0;
 wire n_11548_o_0;
 wire n_11549_o_0;
 wire n_11550_o_0;
 wire n_11551_o_0;
 wire n_11552_o_0;
 wire n_11553_o_0;
 wire n_11554_o_0;
 wire n_11555_o_0;
 wire n_11556_o_0;
 wire n_11557_o_0;
 wire n_11558_o_0;
 wire n_11559_o_0;
 wire n_11560_o_0;
 wire n_11561_o_0;
 wire n_11562_o_0;
 wire n_11563_o_0;
 wire n_11564_o_0;
 wire n_11565_o_0;
 wire n_11566_o_0;
 wire n_11567_o_0;
 wire n_11568_o_0;
 wire n_11569_o_0;
 wire n_11570_o_0;
 wire n_11571_o_0;
 wire n_11572_o_0;
 wire n_11573_o_0;
 wire n_11574_o_0;
 wire n_11575_o_0;
 wire n_11576_o_0;
 wire n_11577_o_0;
 wire n_11578_o_0;
 wire n_11579_o_0;
 wire n_11580_o_0;
 wire n_11581_o_0;
 wire n_11582_o_0;
 wire n_11583_o_0;
 wire n_11584_o_0;
 wire n_11585_o_0;
 wire n_11586_o_0;
 wire n_11587_o_0;
 wire n_11588_o_0;
 wire n_11589_o_0;
 wire n_11590_o_0;
 wire n_11591_o_0;
 wire n_11592_o_0;
 wire n_11593_o_0;
 wire n_11594_o_0;
 wire n_11595_o_0;
 wire n_11596_o_0;
 wire n_11597_o_0;
 wire n_11598_o_0;
 wire n_11599_o_0;
 wire n_11600_o_0;
 wire n_11601_o_0;
 wire n_11602_o_0;
 wire n_11603_o_0;
 wire n_11604_o_0;
 wire n_11605_o_0;
 wire n_11606_o_0;
 wire n_11607_o_0;
 wire n_11608_o_0;
 wire n_11609_o_0;
 wire n_11610_o_0;
 wire n_11611_o_0;
 wire n_11612_o_0;
 wire n_11613_o_0;
 wire n_11614_o_0;
 wire n_11615_o_0;
 wire n_11616_o_0;
 wire n_11617_o_0;
 wire n_11618_o_0;
 wire n_11619_o_0;
 wire n_11620_o_0;
 wire n_11621_o_0;
 wire n_11622_o_0;
 wire n_11623_o_0;
 wire n_11624_o_0;
 wire n_11625_o_0;
 wire n_11626_o_0;
 wire n_11627_o_0;
 wire n_11628_o_0;
 wire n_11629_o_0;
 wire n_11630_o_0;
 wire n_11631_o_0;
 wire n_11632_o_0;
 wire n_11633_o_0;
 wire n_11634_o_0;
 wire n_11635_o_0;
 wire n_11636_o_0;
 wire n_11637_o_0;
 wire n_11638_o_0;
 wire n_11639_o_0;
 wire n_11640_o_0;
 wire n_11641_o_0;
 wire n_11642_o_0;
 wire n_11643_o_0;
 wire n_11644_o_0;
 wire n_11645_o_0;
 wire n_11646_o_0;
 wire n_11647_o_0;
 wire n_11648_o_0;
 wire n_11649_o_0;
 wire n_11650_o_0;
 wire n_11651_o_0;
 wire n_11652_o_0;
 wire n_11653_o_0;
 wire n_11654_o_0;
 wire n_11655_o_0;
 wire n_11656_o_0;
 wire n_11657_o_0;
 wire n_11658_o_0;
 wire n_11659_o_0;
 wire n_11660_o_0;
 wire n_11661_o_0;
 wire n_11662_o_0;
 wire n_11663_o_0;
 wire n_11664_o_0;
 wire n_11665_o_0;
 wire n_11666_o_0;
 wire n_11667_o_0;
 wire n_11668_o_0;
 wire n_11669_o_0;
 wire n_11670_o_0;
 wire n_11671_o_0;
 wire n_11672_o_0;
 wire n_11673_o_0;
 wire n_11674_o_0;
 wire n_11674_o_1;
 wire n_11675_o_0;
 wire n_11676_o_0;
 wire n_11677_o_0;
 wire n_11678_o_0;
 wire n_11679_o_0;
 wire n_11680_o_0;
 wire n_11681_o_0;
 wire n_11681_o_1;
 wire n_11682_o_0;
 wire n_11683_o_0;
 wire n_11684_o_0;
 wire n_11685_o_0;
 wire n_11686_o_0;
 wire n_11687_o_0;
 wire n_11688_o_0;
 wire n_11689_o_0;
 wire n_11690_o_0;
 wire n_11691_o_0;
 wire n_11692_o_0;
 wire n_11693_o_0;
 wire n_11694_o_0;
 wire n_11695_o_0;
 wire n_11696_o_0;
 wire n_11697_o_0;
 wire n_11698_o_0;
 wire n_11699_o_0;
 wire n_11700_o_0;
 wire n_11701_o_0;
 wire n_11702_o_0;
 wire n_11703_o_0;
 wire n_11704_o_0;
 wire n_11705_o_0;
 wire n_11706_o_0;
 wire n_11707_o_0;
 wire n_11708_o_0;
 wire n_11709_o_0;
 wire n_11710_o_0;
 wire n_11711_o_0;
 wire n_11712_o_0;
 wire n_11713_o_0;
 wire n_11714_o_0;
 wire n_11715_o_0;
 wire n_11716_o_0;
 wire n_11717_o_0;
 wire n_11718_o_0;
 wire n_11719_o_0;
 wire n_11720_o_0;
 wire n_11721_o_0;
 wire n_11722_o_0;
 wire n_11723_o_0;
 wire n_11724_o_0;
 wire n_11725_o_0;
 wire n_11726_o_0;
 wire n_11727_o_0;
 wire n_11728_o_0;
 wire n_11729_o_0;
 wire n_11730_o_0;
 wire n_11731_o_0;
 wire n_11732_o_0;
 wire n_11733_o_0;
 wire n_11734_o_0;
 wire n_11735_o_0;
 wire n_11736_o_0;
 wire n_11737_o_0;
 wire n_11738_o_0;
 wire n_11739_o_0;
 wire n_11740_o_0;
 wire n_11741_o_0;
 wire n_11742_o_0;
 wire n_11743_o_0;
 wire n_11744_o_0;
 wire n_11745_o_0;
 wire n_11746_o_0;
 wire n_11747_o_0;
 wire n_11748_o_0;
 wire n_11749_o_0;
 wire n_11749_o_1;
 wire n_11750_o_0;
 wire n_11751_o_0;
 wire n_11752_o_0;
 wire n_11753_o_0;
 wire n_11754_o_0;
 wire n_11755_o_0;
 wire n_11756_o_0;
 wire n_11757_o_0;
 wire n_11758_o_0;
 wire n_11759_o_0;
 wire n_11760_o_0;
 wire n_11761_o_0;
 wire n_11762_o_0;
 wire n_11763_o_0;
 wire n_11764_o_0;
 wire n_11765_o_0;
 wire n_11766_o_0;
 wire n_11767_o_0;
 wire n_11768_o_0;
 wire n_11769_o_0;
 wire n_11770_o_0;
 wire n_11771_o_0;
 wire n_11772_o_0;
 wire n_11773_o_0;
 wire n_11774_o_0;
 wire n_11775_o_0;
 wire n_11776_o_0;
 wire n_11777_o_0;
 wire n_11778_o_0;
 wire n_11779_o_0;
 wire n_11780_o_0;
 wire n_11781_o_0;
 wire n_11782_o_0;
 wire n_11783_o_0;
 wire n_11784_o_0;
 wire n_11785_o_0;
 wire n_11786_o_0;
 wire n_11787_o_0;
 wire n_11788_o_0;
 wire n_11789_o_0;
 wire n_11790_o_0;
 wire n_11791_o_0;
 wire n_11792_o_0;
 wire n_11793_o_0;
 wire n_11794_o_0;
 wire n_11795_o_0;
 wire n_11796_o_0;
 wire n_11797_o_0;
 wire n_11798_o_0;
 wire n_11799_o_0;
 wire n_11800_o_0;
 wire n_11801_o_0;
 wire n_11802_o_0;
 wire n_11803_o_0;
 wire n_11804_o_0;
 wire n_11805_o_0;
 wire n_11806_o_0;
 wire n_11807_o_0;
 wire n_11808_o_0;
 wire n_11809_o_0;
 wire n_11810_o_0;
 wire n_11811_o_0;
 wire n_11812_o_0;
 wire n_11813_o_0;
 wire n_11814_o_0;
 wire n_11815_o_0;
 wire n_11816_o_0;
 wire n_11817_o_0;
 wire n_11818_o_0;
 wire n_11819_o_0;
 wire n_11820_o_0;
 wire n_11821_o_0;
 wire n_11822_o_0;
 wire n_11823_o_0;
 wire n_11824_o_0;
 wire n_11825_o_0;
 wire n_11826_o_0;
 wire n_11827_o_0;
 wire n_11828_o_0;
 wire n_11829_o_0;
 wire n_11830_o_0;
 wire n_11831_o_0;
 wire n_11832_o_0;
 wire n_11833_o_0;
 wire n_11834_o_0;
 wire n_11835_o_0;
 wire n_11836_o_0;
 wire n_11837_o_0;
 wire n_11838_o_0;
 wire n_11839_o_0;
 wire n_11840_o_0;
 wire n_11841_o_0;
 wire n_11842_o_0;
 wire n_11843_o_0;
 wire n_11844_o_0;
 wire n_11845_o_0;
 wire n_11846_o_0;
 wire n_11847_o_0;
 wire n_11848_o_0;
 wire n_11849_o_0;
 wire n_11850_o_0;
 wire n_11851_o_0;
 wire n_11852_o_0;
 wire n_11853_o_0;
 wire n_11854_o_0;
 wire n_11855_o_0;
 wire n_11856_o_0;
 wire n_11857_o_0;
 wire n_11858_o_0;
 wire n_11859_o_0;
 wire n_11860_o_0;
 wire n_11861_o_0;
 wire n_11862_o_0;
 wire n_11863_o_0;
 wire n_11864_o_0;
 wire n_11865_o_0;
 wire n_11866_o_0;
 wire n_11867_o_0;
 wire n_11868_o_0;
 wire n_11869_o_0;
 wire n_11870_o_0;
 wire n_11871_o_0;
 wire n_11872_o_0;
 wire n_11873_o_0;
 wire n_11874_o_0;
 wire n_11875_o_0;
 wire n_11876_o_0;
 wire n_11877_o_0;
 wire n_11878_o_0;
 wire n_11879_o_0;
 wire n_11880_o_0;
 wire n_11881_o_0;
 wire n_11882_o_0;
 wire n_11883_o_0;
 wire n_11884_o_0;
 wire n_11885_o_0;
 wire n_11886_o_0;
 wire n_11887_o_0;
 wire n_11888_o_0;
 wire n_11889_o_0;
 wire n_11890_o_0;
 wire n_11891_o_0;
 wire n_11892_o_0;
 wire n_11893_o_0;
 wire n_11894_o_0;
 wire n_11895_o_0;
 wire n_11896_o_0;
 wire n_11897_o_0;
 wire n_11898_o_0;
 wire n_11899_o_0;
 wire n_11900_o_0;
 wire n_11901_o_0;
 wire n_11902_o_0;
 wire n_11903_o_0;
 wire n_11904_o_0;
 wire n_11905_o_0;
 wire n_11906_o_0;
 wire n_11907_o_0;
 wire n_11908_o_0;
 wire n_11909_o_0;
 wire n_11910_o_0;
 wire n_11911_o_0;
 wire n_11912_o_0;
 wire n_11913_o_0;
 wire n_11914_o_0;
 wire n_11915_o_0;
 wire n_11916_o_0;
 wire n_11917_o_0;
 wire n_11918_o_0;
 wire n_11919_o_0;
 wire n_11920_o_0;
 wire n_11921_o_0;
 wire n_11922_o_0;
 wire n_11923_o_0;
 wire n_11924_o_0;
 wire n_11925_o_0;
 wire n_11926_o_0;
 wire n_11927_o_0;
 wire n_11928_o_0;
 wire n_11929_o_0;
 wire n_11930_o_0;
 wire n_11931_o_0;
 wire n_11932_o_0;
 wire n_11933_o_0;
 wire n_11934_o_0;
 wire n_11935_o_0;
 wire n_11936_o_0;
 wire n_11937_o_0;
 wire n_11938_o_0;
 wire n_11939_o_0;
 wire n_11940_o_0;
 wire n_11941_o_0;
 wire n_11942_o_0;
 wire n_11943_o_0;
 wire n_11944_o_0;
 wire n_11945_o_0;
 wire n_11946_o_0;
 wire n_11947_o_0;
 wire n_11948_o_0;
 wire n_11949_o_0;
 wire n_11950_o_0;
 wire n_11951_o_0;
 wire n_11952_o_0;
 wire n_11953_o_0;
 wire n_11954_o_0;
 wire n_11955_o_0;
 wire n_11956_o_0;
 wire n_11957_o_0;
 wire n_11958_o_0;
 wire n_11959_o_0;
 wire n_11960_o_0;
 wire n_11961_o_0;
 wire n_11962_o_0;
 wire n_11963_o_0;
 wire n_11964_o_0;
 wire n_11965_o_0;
 wire n_11966_o_0;
 wire n_11967_o_0;
 wire n_11968_o_0;
 wire n_11969_o_0;
 wire n_11970_o_0;
 wire n_11971_o_0;
 wire n_11972_o_0;
 wire n_11973_o_0;
 wire n_11974_o_0;
 wire n_11975_o_0;
 wire n_11976_o_0;
 wire n_11977_o_0;
 wire n_11978_o_0;
 wire n_11979_o_0;
 wire n_11980_o_0;
 wire n_11981_o_0;
 wire n_11982_o_0;
 wire n_11983_o_0;
 wire n_11984_o_0;
 wire n_11985_o_0;
 wire n_11986_o_0;
 wire n_11987_o_0;
 wire n_11988_o_0;
 wire n_11989_o_0;
 wire n_11990_o_0;
 wire n_11991_o_0;
 wire n_11992_o_0;
 wire n_11993_o_0;
 wire n_11994_o_0;
 wire n_11995_o_0;
 wire n_11996_o_0;
 wire n_11997_o_0;
 wire n_11998_o_0;
 wire n_11999_o_0;
 wire n_12000_o_0;
 wire n_12001_o_0;
 wire n_12002_o_0;
 wire n_12003_o_0;
 wire n_12004_o_0;
 wire n_12005_o_0;
 wire n_12006_o_0;
 wire n_12007_o_0;
 wire n_12008_o_0;
 wire n_12009_o_0;
 wire n_12010_o_0;
 wire n_12011_o_0;
 wire n_12012_o_0;
 wire n_12013_o_0;
 wire n_12014_o_0;
 wire n_12015_o_0;
 wire n_12016_o_0;
 wire n_12017_o_0;
 wire n_12018_o_0;
 wire n_12019_o_0;
 wire n_12020_o_0;
 wire n_12021_o_0;
 wire n_12022_o_0;
 wire n_12023_o_0;
 wire n_12024_o_0;
 wire n_12025_o_0;
 wire n_12026_o_0;
 wire n_12027_o_0;
 wire n_12028_o_0;
 wire n_12029_o_0;
 wire n_12030_o_0;
 wire n_12031_o_0;
 wire n_12032_o_0;
 wire n_12033_o_0;
 wire n_12034_o_0;
 wire n_12035_o_0;
 wire n_12036_o_0;
 wire n_12037_o_0;
 wire n_12038_o_0;
 wire n_12039_o_0;
 wire n_12040_o_0;
 wire n_12041_o_0;
 wire n_12042_o_0;
 wire n_12043_o_0;
 wire n_12044_o_0;
 wire n_12045_o_0;
 wire n_12046_o_0;
 wire n_12047_o_0;
 wire n_12048_o_0;
 wire n_12049_o_0;
 wire n_12050_o_0;
 wire n_12051_o_0;
 wire n_12052_o_0;
 wire n_12053_o_0;
 wire n_12054_o_0;
 wire n_12055_o_0;
 wire n_12056_o_0;
 wire n_12057_o_0;
 wire n_12058_o_0;
 wire n_12059_o_0;
 wire n_12060_o_0;
 wire n_12061_o_0;
 wire n_12062_o_0;
 wire n_12063_o_0;
 wire n_12064_o_0;
 wire n_12065_o_0;
 wire n_12066_o_0;
 wire n_12067_o_0;
 wire n_12068_o_0;
 wire n_12069_o_0;
 wire n_12070_o_0;
 wire n_12071_o_0;
 wire n_12072_o_0;
 wire n_12073_o_0;
 wire n_12074_o_0;
 wire n_12075_o_0;
 wire n_12076_o_0;
 wire n_12077_o_0;
 wire n_12078_o_0;
 wire n_12079_o_0;
 wire n_12080_o_0;
 wire n_12081_o_0;
 wire n_12082_o_0;
 wire n_12083_o_0;
 wire n_12084_o_0;
 wire n_12085_o_0;
 wire n_12086_o_0;
 wire n_12087_o_0;
 wire n_12088_o_0;
 wire n_12089_o_0;
 wire n_12090_o_0;
 wire n_12091_o_0;
 wire n_12092_o_0;
 wire n_12093_o_0;
 wire n_12094_o_0;
 wire n_12095_o_0;
 wire n_12096_o_0;
 wire n_12097_o_0;
 wire n_12098_o_0;
 wire n_12099_o_0;
 wire n_12100_o_0;
 wire n_12101_o_0;
 wire n_12102_o_0;
 wire n_12103_o_0;
 wire n_12104_o_0;
 wire n_12105_o_0;
 wire n_12106_o_0;
 wire n_12107_o_0;
 wire n_12108_o_0;
 wire n_12109_o_0;
 wire n_12110_o_0;
 wire n_12111_o_0;
 wire n_12112_o_0;
 wire n_12113_o_0;
 wire n_12114_o_0;
 wire n_12115_o_0;
 wire n_12116_o_0;
 wire n_12117_o_0;
 wire n_12118_o_0;
 wire n_12119_o_0;
 wire n_12120_o_0;
 wire n_12121_o_0;
 wire n_12122_o_0;
 wire n_12123_o_0;
 wire n_12124_o_0;
 wire n_12125_o_0;
 wire n_12126_o_0;
 wire n_12127_o_0;
 wire n_12128_o_0;
 wire n_12129_o_0;
 wire n_12130_o_0;
 wire n_12131_o_0;
 wire n_12132_o_0;
 wire n_12133_o_0;
 wire n_12134_o_0;
 wire n_12135_o_0;
 wire n_12136_o_0;
 wire n_12137_o_0;
 wire n_12138_o_0;
 wire n_12139_o_0;
 wire n_12140_o_0;
 wire n_12141_o_0;
 wire n_12142_o_0;
 wire n_12143_o_0;
 wire n_12144_o_0;
 wire n_12145_o_0;
 wire n_12146_o_0;
 wire n_12147_o_0;
 wire n_12148_o_0;
 wire n_12149_o_0;
 wire n_12150_o_0;
 wire n_12151_o_0;
 wire n_12152_o_0;
 wire n_12153_o_0;
 wire n_12154_o_0;
 wire n_12155_o_0;
 wire n_12156_o_0;
 wire n_12157_o_0;
 wire n_12158_o_0;
 wire n_12159_o_0;
 wire n_12160_o_0;
 wire n_12161_o_0;
 wire n_12162_o_0;
 wire n_12163_o_0;
 wire n_12164_o_0;
 wire n_12165_o_0;
 wire n_12166_o_0;
 wire n_12167_o_0;
 wire n_12168_o_0;
 wire n_12169_o_0;
 wire n_12170_o_0;
 wire n_12171_o_0;
 wire n_12172_o_0;
 wire n_12173_o_0;
 wire n_12174_o_0;
 wire n_12175_o_0;
 wire n_12176_o_0;
 wire n_12177_o_0;
 wire n_12178_o_0;
 wire n_12179_o_0;
 wire n_12180_o_0;
 wire n_12181_o_0;
 wire n_12182_o_0;
 wire n_12183_o_0;
 wire n_12184_o_0;
 wire n_12185_o_0;
 wire n_12186_o_0;
 wire n_12187_o_0;
 wire n_12188_o_0;
 wire n_12189_o_0;
 wire n_12190_o_0;
 wire n_12191_o_0;
 wire n_12192_o_0;
 wire n_12193_o_0;
 wire n_12194_o_0;
 wire n_12195_o_0;
 wire n_12196_o_0;
 wire n_12197_o_0;
 wire n_12198_o_0;
 wire n_12199_o_0;
 wire n_12200_o_0;
 wire n_12201_o_0;
 wire n_12202_o_0;
 wire n_12203_o_0;
 wire n_12204_o_0;
 wire n_12205_o_0;
 wire n_12206_o_0;
 wire n_12207_o_0;
 wire n_12208_o_0;
 wire n_12209_o_0;
 wire n_12210_o_0;
 wire n_12211_o_0;
 wire n_12212_o_0;
 wire n_12213_o_0;
 wire n_12214_o_0;
 wire n_12215_o_0;
 wire n_12216_o_0;
 wire n_12217_o_0;
 wire n_12218_o_0;
 wire n_12219_o_0;
 wire n_12220_o_0;
 wire n_12221_o_0;
 wire n_12222_o_0;
 wire n_12223_o_0;
 wire n_12224_o_0;
 wire n_12225_o_0;
 wire n_12226_o_0;
 wire n_12227_o_0;
 wire n_12228_o_0;
 wire n_12229_o_0;
 wire n_12230_o_0;
 wire n_12231_o_0;
 wire n_12232_o_0;
 wire n_12233_o_0;
 wire n_12234_o_0;
 wire n_12235_o_0;
 wire n_12236_o_0;
 wire n_12237_o_0;
 wire n_12238_o_0;
 wire n_12239_o_0;
 wire n_12240_o_0;
 wire n_12241_o_0;
 wire n_12242_o_0;
 wire n_12243_o_0;
 wire n_12244_o_0;
 wire n_12245_o_0;
 wire n_12246_o_0;
 wire n_12247_o_0;
 wire n_12248_o_0;
 wire n_12249_o_0;
 wire n_12250_o_0;
 wire n_12251_o_0;
 wire n_12252_o_0;
 wire n_12253_o_0;
 wire n_12254_o_0;
 wire n_12255_o_0;
 wire n_12256_o_0;
 wire n_12257_o_0;
 wire n_12258_o_0;
 wire n_12259_o_0;
 wire n_12260_o_0;
 wire n_12261_o_0;
 wire n_12262_o_0;
 wire n_12263_o_0;
 wire n_12264_o_0;
 wire n_12265_o_0;
 wire n_12266_o_0;
 wire n_12267_o_0;
 wire n_12268_o_0;
 wire n_12269_o_0;
 wire n_12270_o_0;
 wire n_12271_o_0;
 wire n_12272_o_0;
 wire n_12273_o_0;
 wire n_12274_o_0;
 wire n_12275_o_0;
 wire n_12276_o_0;
 wire n_12277_o_0;
 wire n_12278_o_0;
 wire n_12279_o_0;
 wire n_12280_o_0;
 wire n_12281_o_0;
 wire n_12282_o_0;
 wire n_12283_o_0;
 wire n_12284_o_0;
 wire n_12285_o_0;
 wire n_12286_o_0;
 wire n_12287_o_0;
 wire n_12288_o_0;
 wire n_12289_o_0;
 wire n_12290_o_0;
 wire n_12291_o_0;
 wire n_12292_o_0;
 wire n_12293_o_0;
 wire n_12294_o_0;
 wire n_12295_o_0;
 wire n_12296_o_0;
 wire n_12297_o_0;
 wire n_12298_o_0;
 wire n_12299_o_0;
 wire n_12300_o_0;
 wire n_12301_o_0;
 wire n_12302_o_0;
 wire n_12303_o_0;
 wire n_12304_o_0;
 wire n_12305_o_0;
 wire n_12306_o_0;
 wire n_12307_o_0;
 wire n_12308_o_0;
 wire n_12309_o_0;
 wire n_12310_o_0;
 wire n_12311_o_0;
 wire n_12312_o_0;
 wire n_12313_o_0;
 wire n_12314_o_0;
 wire n_12315_o_0;
 wire n_12316_o_0;
 wire n_12317_o_0;
 wire n_12318_o_0;
 wire n_12319_o_0;
 wire n_12320_o_0;
 wire n_12321_o_0;
 wire n_12322_o_0;
 wire n_12323_o_0;
 wire n_12324_o_0;
 wire n_12325_o_0;
 wire n_12326_o_0;
 wire n_12327_o_0;
 wire n_12328_o_0;
 wire n_12329_o_0;
 wire n_12330_o_0;
 wire n_12331_o_0;
 wire n_12332_o_0;
 wire n_12333_o_0;
 wire n_12334_o_0;
 wire n_12335_o_0;
 wire n_12336_o_0;
 wire n_12337_o_0;
 wire n_12338_o_0;
 wire n_12339_o_0;
 wire n_12340_o_0;
 wire n_12341_o_0;
 wire n_12342_o_0;
 wire n_12343_o_0;
 wire n_12344_o_0;
 wire n_12345_o_0;
 wire n_12346_o_0;
 wire n_12347_o_0;
 wire n_12348_o_0;
 wire n_12349_o_0;
 wire n_12350_o_0;
 wire n_12351_o_0;
 wire n_12352_o_0;
 wire n_12353_o_0;
 wire n_12354_o_0;
 wire n_12355_o_0;
 wire n_12356_o_0;
 wire n_12357_o_0;
 wire n_12358_o_0;
 wire n_12359_o_0;
 wire n_12360_o_0;
 wire n_12361_o_0;
 wire n_12362_o_0;
 wire n_12363_o_0;
 wire n_12364_o_0;
 wire n_12365_o_0;
 wire n_12366_o_0;
 wire n_12367_o_0;
 wire n_12368_o_0;
 wire n_12369_o_0;
 wire n_12370_o_0;
 wire n_12371_o_0;
 wire n_12372_o_0;
 wire n_12373_o_0;
 wire n_12374_o_0;
 wire n_12375_o_0;
 wire n_12376_o_0;
 wire n_12377_o_0;
 wire n_12378_o_0;
 wire n_12379_o_0;
 wire n_12380_o_0;
 wire n_12381_o_0;
 wire n_12382_o_0;
 wire n_12383_o_0;
 wire n_12384_o_0;
 wire n_12385_o_0;
 wire n_12386_o_0;
 wire n_12387_o_0;
 wire n_12388_o_0;
 wire n_12389_o_0;
 wire n_12390_o_0;
 wire n_12391_o_0;
 wire n_12392_o_0;
 wire n_12393_o_0;
 wire n_12394_o_0;
 wire n_12395_o_0;
 wire n_12396_o_0;
 wire n_12397_o_0;
 wire n_12398_o_0;
 wire n_12399_o_0;
 wire n_12400_o_0;
 wire n_12401_o_0;
 wire n_12402_o_0;
 wire n_12403_o_0;
 wire n_12404_o_0;
 wire n_12405_o_0;
 wire n_12406_o_0;
 wire n_12407_o_0;
 wire n_12408_o_0;
 wire n_12409_o_0;
 wire n_12410_o_0;
 wire n_12411_o_0;
 wire n_12412_o_0;
 wire n_12413_o_0;
 wire n_12414_o_0;
 wire n_12415_o_0;
 wire n_12416_o_0;
 wire n_12417_o_0;
 wire n_12418_o_0;
 wire n_12419_o_0;
 wire n_12420_o_0;
 wire n_12421_o_0;
 wire n_12422_o_0;
 wire n_12423_o_0;
 wire n_12424_o_0;
 wire n_12425_o_0;
 wire n_12426_o_0;
 wire n_12427_o_0;
 wire n_12428_o_0;
 wire n_12429_o_0;
 wire n_12430_o_0;
 wire n_12431_o_0;
 wire n_12432_o_0;
 wire n_12433_o_0;
 wire n_12434_o_0;
 wire n_12435_o_0;
 wire n_12436_o_0;
 wire n_12437_o_0;
 wire n_12438_o_0;
 wire n_12439_o_0;
 wire n_12440_o_0;
 wire n_12441_o_0;
 wire n_12442_o_0;
 wire n_12443_o_0;
 wire n_12444_o_0;
 wire n_12445_o_0;
 wire n_12446_o_0;
 wire n_12447_o_0;
 wire n_12448_o_0;
 wire n_12449_o_0;
 wire n_12450_o_0;
 wire n_12451_o_0;
 wire n_12452_o_0;
 wire n_12453_o_0;
 wire n_12454_o_0;
 wire n_12455_o_0;
 wire n_12456_o_0;
 wire n_12457_o_0;
 wire n_12458_o_0;
 wire n_12459_o_0;
 wire n_12460_o_0;
 wire n_12461_o_0;
 wire n_12462_o_0;
 wire n_12463_o_0;
 wire n_12464_o_0;
 wire n_12465_o_0;
 wire n_12466_o_0;
 wire n_12467_o_0;
 wire n_12468_o_0;
 wire n_12469_o_0;
 wire n_12470_o_0;
 wire n_12471_o_0;
 wire n_12472_o_0;
 wire n_12473_o_0;
 wire n_12474_o_0;
 wire n_12475_o_0;
 wire n_12476_o_0;
 wire n_12477_o_0;
 wire n_12478_o_0;
 wire n_12479_o_0;
 wire n_12480_o_0;
 wire n_12481_o_0;
 wire n_12482_o_0;
 wire n_12483_o_0;
 wire n_12484_o_0;
 wire n_12485_o_0;
 wire n_12486_o_0;
 wire n_12487_o_0;
 wire n_12488_o_0;
 wire n_12489_o_0;
 wire n_12490_o_0;
 wire n_12491_o_0;
 wire n_12492_o_0;
 wire n_12493_o_0;
 wire n_12494_o_0;
 wire n_12495_o_0;
 wire n_12496_o_0;
 wire n_12497_o_0;
 wire n_12498_o_0;
 wire n_12499_o_0;
 wire n_12500_o_0;
 wire n_12501_o_0;
 wire n_12502_o_0;
 wire n_12503_o_0;
 wire n_12504_o_0;
 wire n_12505_o_0;
 wire n_12506_o_0;
 wire n_12507_o_0;
 wire n_12508_o_0;
 wire n_12509_o_0;
 wire n_12510_o_0;
 wire n_12511_o_0;
 wire n_12512_o_0;
 wire n_12513_o_0;
 wire n_12514_o_0;
 wire n_12515_o_0;
 wire n_12516_o_0;
 wire n_12517_o_0;
 wire n_12518_o_0;
 wire n_12519_o_0;
 wire n_12520_o_0;
 wire n_12521_o_0;
 wire n_12522_o_0;
 wire n_12523_o_0;
 wire n_12524_o_0;
 wire n_12525_o_0;
 wire n_12526_o_0;
 wire n_12527_o_0;
 wire n_12528_o_0;
 wire n_12529_o_0;
 wire n_12530_o_0;
 wire n_12531_o_0;
 wire n_12532_o_0;
 wire n_12533_o_0;
 wire n_12534_o_0;
 wire n_12535_o_0;
 wire n_12536_o_0;
 wire n_12537_o_0;
 wire n_12538_o_0;
 wire n_12539_o_0;
 wire n_12540_o_0;
 wire n_12541_o_0;
 wire n_12542_o_0;
 wire n_12543_o_0;
 wire n_12544_o_0;
 wire n_12545_o_0;
 wire n_12546_o_0;
 wire n_12547_o_0;
 wire n_12548_o_0;
 wire n_12549_o_0;
 wire n_12550_o_0;
 wire n_12551_o_0;
 wire n_12552_o_0;
 wire n_12553_o_0;
 wire n_12554_o_0;
 wire n_12555_o_0;
 wire n_12556_o_0;
 wire n_12557_o_0;
 wire n_12558_o_0;
 wire n_12559_o_0;
 wire n_12560_o_0;
 wire n_12561_o_0;
 wire n_12562_o_0;
 wire n_12563_o_0;
 wire n_12564_o_0;
 wire n_12565_o_0;
 wire n_12566_o_0;
 wire n_12567_o_0;
 wire n_12568_o_0;
 wire n_12569_o_0;
 wire n_12570_o_0;
 wire n_12571_o_0;
 wire n_12572_o_0;
 wire n_12573_o_0;
 wire n_12574_o_0;
 wire n_12575_o_0;
 wire n_12576_o_0;
 wire n_12577_o_0;
 wire n_12578_o_0;
 wire n_12579_o_0;
 wire n_12580_o_0;
 wire n_12581_o_0;
 wire n_12582_o_0;
 wire n_12583_o_0;
 wire n_12584_o_0;
 wire n_12585_o_0;
 wire n_12586_o_0;
 wire n_12587_o_0;
 wire n_12588_o_0;
 wire n_12589_o_0;
 wire n_12590_o_0;
 wire n_12591_o_0;
 wire n_12592_o_0;
 wire n_12593_o_0;
 wire n_12594_o_0;
 wire n_12595_o_0;
 wire n_12596_o_0;
 wire n_12597_o_0;
 wire n_12598_o_0;
 wire n_12599_o_0;
 wire n_12600_o_0;
 wire n_12601_o_0;
 wire n_12602_o_0;
 wire n_12603_o_0;
 wire n_12604_o_0;
 wire n_12605_o_0;
 wire n_12606_o_0;
 wire n_12607_o_0;
 wire n_12608_o_0;
 wire n_12609_o_0;
 wire n_12610_o_0;
 wire n_12611_o_0;
 wire n_12612_o_0;
 wire n_12613_o_0;
 wire n_12614_o_0;
 wire n_12615_o_0;
 wire n_12616_o_0;
 wire n_12617_o_0;
 wire n_12618_o_0;
 wire n_12619_o_0;
 wire n_12620_o_0;
 wire n_12621_o_0;
 wire n_12622_o_0;
 wire n_12623_o_0;
 wire n_12624_o_0;
 wire n_12625_o_0;
 wire n_12626_o_0;
 wire n_12627_o_0;
 wire n_12628_o_0;
 wire n_12629_o_0;
 wire n_12630_o_0;
 wire n_12631_o_0;
 wire n_12632_o_0;
 wire n_12633_o_0;
 wire n_12634_o_0;
 wire n_12635_o_0;
 wire n_12636_o_0;
 wire n_12637_o_0;
 wire n_12638_o_0;
 wire n_12639_o_0;
 wire n_12640_o_0;
 wire n_12641_o_0;
 wire n_12642_o_0;
 wire n_12643_o_0;
 wire n_12644_o_0;
 wire n_12645_o_0;
 wire n_12646_o_0;
 wire n_12647_o_0;
 wire n_12648_o_0;
 wire n_12649_o_0;
 wire n_12650_o_0;
 wire n_12651_o_0;
 wire n_12652_o_0;
 wire n_12653_o_0;
 wire n_12654_o_0;
 wire n_12655_o_0;
 wire n_12656_o_0;
 wire n_12657_o_0;
 wire n_12658_o_0;
 wire n_12659_o_0;
 wire n_12660_o_0;
 wire n_12661_o_0;
 wire n_12662_o_0;
 wire n_12663_o_0;
 wire n_12664_o_0;
 wire n_12665_o_0;
 wire n_12666_o_0;
 wire n_12667_o_0;
 wire n_12668_o_0;
 wire n_12669_o_0;
 wire n_12670_o_0;
 wire n_12671_o_0;
 wire n_12672_o_0;
 wire n_12673_o_0;
 wire n_12674_o_0;
 wire n_12675_o_0;
 wire n_12676_o_0;
 wire n_12677_o_0;
 wire n_12678_o_0;
 wire n_12679_o_0;
 wire n_12680_o_0;
 wire n_12681_o_0;
 wire n_12682_o_0;
 wire n_12683_o_0;
 wire n_12684_o_0;
 wire n_12685_o_0;
 wire n_12686_o_0;
 wire n_12687_o_0;
 wire n_12688_o_0;
 wire n_12689_o_0;
 wire n_12690_o_0;
 wire n_12691_o_0;
 wire n_12692_o_0;
 wire n_12693_o_0;
 wire n_12694_o_0;
 wire n_12695_o_0;
 wire n_12696_o_0;
 wire n_12697_o_0;
 wire n_12698_o_0;
 wire n_12699_o_0;
 wire n_12700_o_0;
 wire n_12701_o_0;
 wire n_12702_o_0;
 wire n_12703_o_0;
 wire n_12704_o_0;
 wire n_12705_o_0;
 wire n_12706_o_0;
 wire n_12707_o_0;
 wire n_12708_o_0;
 wire n_12709_o_0;
 wire n_12710_o_0;
 wire n_12711_o_0;
 wire n_12712_o_0;
 wire n_12713_o_0;
 wire n_12714_o_0;
 wire n_12715_o_0;
 wire n_12716_o_0;
 wire n_12717_o_0;
 wire n_12718_o_0;
 wire n_12719_o_0;
 wire n_12720_o_0;
 wire n_12721_o_0;
 wire n_12722_o_0;
 wire n_12723_o_0;
 wire n_12724_o_0;
 wire n_12725_o_0;
 wire n_12726_o_0;
 wire n_12727_o_0;
 wire n_12728_o_0;
 wire n_12729_o_0;
 wire n_12730_o_0;
 wire n_12731_o_0;
 wire n_12732_o_0;
 wire n_12733_o_0;
 wire n_12734_o_0;
 wire n_12735_o_0;
 wire n_12736_o_0;
 wire n_12737_o_0;
 wire n_12738_o_0;
 wire n_12739_o_0;
 wire n_12740_o_0;
 wire n_12741_o_0;
 wire n_12742_o_0;
 wire n_12743_o_0;
 wire n_12744_o_0;
 wire n_12745_o_0;
 wire n_12746_o_0;
 wire n_12747_o_0;
 wire n_12748_o_0;
 wire n_12749_o_0;
 wire n_12750_o_0;
 wire n_12751_o_0;
 wire n_12752_o_0;
 wire n_12753_o_0;
 wire n_12754_o_0;
 wire n_12755_o_0;
 wire n_12756_o_0;
 wire n_12757_o_0;
 wire n_12758_o_0;
 wire n_12759_o_0;
 wire n_12760_o_0;
 wire n_12761_o_0;
 wire n_12762_o_0;
 wire n_12763_o_0;
 wire n_12764_o_0;
 wire n_12765_o_0;
 wire n_12766_o_0;
 wire n_12767_o_0;
 wire n_12768_o_0;
 wire n_12769_o_0;
 wire n_12770_o_0;
 wire n_12771_o_0;
 wire n_12772_o_0;
 wire n_12773_o_0;
 wire n_12774_o_0;
 wire n_12775_o_0;
 wire n_12776_o_0;
 wire n_12777_o_0;
 wire n_12778_o_0;
 wire n_12779_o_0;
 wire n_12780_o_0;
 wire n_12781_o_0;
 wire n_12782_o_0;
 wire n_12783_o_0;
 wire n_12784_o_0;
 wire n_12785_o_0;
 wire n_12786_o_0;
 wire n_12787_o_0;
 wire n_12788_o_0;
 wire n_12789_o_0;
 wire n_12790_o_0;
 wire n_12791_o_0;
 wire n_12792_o_0;
 wire n_12793_o_0;
 wire n_12794_o_0;
 wire n_12795_o_0;
 wire n_12796_o_0;
 wire n_12797_o_0;
 wire n_12798_o_0;
 wire n_12799_o_0;
 wire n_12800_o_0;
 wire n_12801_o_0;
 wire n_12802_o_0;
 wire n_12803_o_0;
 wire n_12804_o_0;
 wire n_12805_o_0;
 wire n_12806_o_0;
 wire n_12807_o_0;
 wire n_12808_o_0;
 wire n_12809_o_0;
 wire n_12810_o_0;
 wire n_12811_o_0;
 wire n_12812_o_0;
 wire n_12813_o_0;
 wire n_12814_o_0;
 wire n_12815_o_0;
 wire n_12816_o_0;
 wire n_12817_o_0;
 wire n_12818_o_0;
 wire n_12819_o_0;
 wire n_12820_o_0;
 wire n_12821_o_0;
 wire n_12822_o_0;
 wire n_12823_o_0;
 wire n_12824_o_0;
 wire n_12825_o_0;
 wire n_12826_o_0;
 wire n_12827_o_0;
 wire n_12828_o_0;
 wire n_12829_o_0;
 wire n_12830_o_0;
 wire n_12831_o_0;
 wire n_12832_o_0;
 wire n_12833_o_0;
 wire n_12834_o_0;
 wire n_12835_o_0;
 wire n_12836_o_0;
 wire n_12837_o_0;
 wire n_12838_o_0;
 wire n_12839_o_0;
 wire n_12840_o_0;
 wire n_12841_o_0;
 wire n_12842_o_0;
 wire n_12843_o_0;
 wire n_12844_o_0;
 wire n_12845_o_0;
 wire n_12846_o_0;
 wire n_12847_o_0;
 wire n_12848_o_0;
 wire n_12849_o_0;
 wire n_12850_o_0;
 wire n_12851_o_0;
 wire n_12852_o_0;
 wire n_12853_o_0;
 wire n_12854_o_0;
 wire n_12855_o_0;
 wire n_12856_o_0;
 wire n_12857_o_0;
 wire n_12858_o_0;
 wire n_12859_o_0;
 wire n_12860_o_0;
 wire n_12861_o_0;
 wire n_12862_o_0;
 wire n_12863_o_0;
 wire n_12864_o_0;
 wire n_12865_o_0;
 wire n_12866_o_0;
 wire n_12867_o_0;
 wire n_12868_o_0;
 wire n_12869_o_0;
 wire n_12870_o_0;
 wire n_12871_o_0;
 wire n_12872_o_0;
 wire n_12873_o_0;
 wire n_12874_o_0;
 wire n_12875_o_0;
 wire n_12876_o_0;
 wire n_12877_o_0;
 wire n_12878_o_0;
 wire n_12879_o_0;
 wire n_12880_o_0;
 wire n_12881_o_0;
 wire n_12882_o_0;
 wire n_12883_o_0;
 wire n_12884_o_0;
 wire n_12885_o_0;
 wire n_12886_o_0;
 wire n_12887_o_0;
 wire n_12888_o_0;
 wire n_12889_o_0;
 wire n_12890_o_0;
 wire n_12891_o_0;
 wire n_12892_o_0;
 wire n_12893_o_0;
 wire n_12894_o_0;
 wire n_12895_o_0;
 wire n_12896_o_0;
 wire n_12897_o_0;
 wire n_12898_o_0;
 wire n_12899_o_0;
 wire n_12900_o_0;
 wire n_12901_o_0;
 wire n_12902_o_0;
 wire n_12903_o_0;
 wire n_12904_o_0;
 wire n_12905_o_0;
 wire n_12906_o_0;
 wire n_12907_o_0;
 wire n_12908_o_0;
 wire n_12909_o_0;
 wire n_12910_o_0;
 wire n_12911_o_0;
 wire n_12912_o_0;
 wire n_12913_o_0;
 wire n_12914_o_0;
 wire n_12915_o_0;
 wire n_12916_o_0;
 wire n_12917_o_0;
 wire n_12918_o_0;
 wire n_12919_o_0;
 wire n_12920_o_0;
 wire n_12921_o_0;
 wire n_12922_o_0;
 wire n_12923_o_0;
 wire n_12924_o_0;
 wire n_12925_o_0;
 wire n_12926_o_0;
 wire n_12927_o_0;
 wire n_12928_o_0;
 wire n_12929_o_0;
 wire n_12930_o_0;
 wire n_12931_o_0;
 wire n_12932_o_0;
 wire n_12933_o_0;
 wire n_12934_o_0;
 wire n_12935_o_0;
 wire n_12936_o_0;
 wire n_12937_o_0;
 wire n_12938_o_0;
 wire n_12939_o_0;
 wire n_12940_o_0;
 wire n_12941_o_0;
 wire n_12942_o_0;
 wire n_12943_o_0;
 wire n_12944_o_0;
 wire n_12945_o_0;
 wire n_12946_o_0;
 wire n_12947_o_0;
 wire n_12948_o_0;
 wire n_12949_o_0;
 wire n_12950_o_0;
 wire n_12951_o_0;
 wire n_12952_o_0;
 wire n_12953_o_0;
 wire n_12954_o_0;
 wire n_12955_o_0;
 wire n_12956_o_0;
 wire n_12957_o_0;
 wire n_12958_o_0;
 wire n_12959_o_0;
 wire n_12960_o_0;
 wire n_12961_o_0;
 wire n_12962_o_0;
 wire n_12963_o_0;
 wire n_12964_o_0;
 wire n_12965_o_0;
 wire n_12966_o_0;
 wire n_12967_o_0;
 wire n_12968_o_0;
 wire n_12969_o_0;
 wire n_12970_o_0;
 wire n_12971_o_0;
 wire n_12972_o_0;
 wire n_12973_o_0;
 wire n_12974_o_0;
 wire n_12975_o_0;
 wire n_12976_o_0;
 wire n_12977_o_0;
 wire n_12978_o_0;
 wire n_12979_o_0;
 wire n_12980_o_0;
 wire n_12981_o_0;
 wire n_12982_o_0;
 wire n_12983_o_0;
 wire n_12984_o_0;
 wire n_12985_o_0;
 wire n_12986_o_0;
 wire n_12987_o_0;
 wire n_12988_o_0;
 wire n_12989_o_0;
 wire n_12990_o_0;
 wire n_12991_o_0;
 wire n_12992_o_0;
 wire n_12993_o_0;
 wire n_12994_o_0;
 wire n_12995_o_0;
 wire n_12996_o_0;
 wire n_12997_o_0;
 wire n_12998_o_0;
 wire n_12999_o_0;
 wire n_13000_o_0;
 wire n_13001_o_0;
 wire n_13002_o_0;
 wire n_13003_o_0;
 wire n_13004_o_0;
 wire n_13005_o_0;
 wire n_13006_o_0;
 wire n_13007_o_0;
 wire n_13008_o_0;
 wire n_13009_o_0;
 wire n_13010_o_0;
 wire n_13011_o_0;
 wire n_13012_o_0;
 wire n_13013_o_0;
 wire n_13014_o_0;
 wire n_13015_o_0;
 wire n_13016_o_0;
 wire n_13017_o_0;
 wire n_13018_o_0;
 wire n_13019_o_0;
 wire n_13020_o_0;
 wire n_13021_o_0;
 wire n_13022_o_0;
 wire n_13023_o_0;
 wire n_13024_o_0;
 wire n_13025_o_0;
 wire n_13026_o_0;
 wire n_13027_o_0;
 wire n_13028_o_0;
 wire n_13029_o_0;
 wire n_13030_o_0;
 wire n_13031_o_0;
 wire n_13032_o_0;
 wire n_13033_o_0;
 wire n_13034_o_0;
 wire n_13035_o_0;
 wire n_13036_o_0;
 wire n_13037_o_0;
 wire n_13038_o_0;
 wire n_13039_o_0;
 wire n_13040_o_0;
 wire n_13041_o_0;
 wire n_13042_o_0;
 wire n_13043_o_0;
 wire n_13044_o_0;
 wire n_13045_o_0;
 wire n_13046_o_0;
 wire n_13047_o_0;
 wire n_13048_o_0;
 wire n_13049_o_0;
 wire n_13050_o_0;
 wire n_13051_o_0;
 wire n_13052_o_0;
 wire n_13053_o_0;
 wire n_13054_o_0;
 wire n_13055_o_0;
 wire n_13056_o_0;
 wire n_13057_o_0;
 wire n_13058_o_0;
 wire n_13059_o_0;
 wire n_13060_o_0;
 wire n_13061_o_0;
 wire n_13062_o_0;
 wire n_13063_o_0;
 wire n_13064_o_0;
 wire n_13065_o_0;
 wire n_13066_o_0;
 wire n_13067_o_0;
 wire n_13068_o_0;
 wire n_13069_o_0;
 wire n_13070_o_0;
 wire n_13071_o_0;
 wire n_13072_o_0;
 wire n_13073_o_0;
 wire n_13074_o_0;
 wire n_13075_o_0;
 wire n_13076_o_0;
 wire n_13077_o_0;
 wire n_13078_o_0;
 wire n_13079_o_0;
 wire n_13080_o_0;
 wire n_13081_o_0;
 wire n_13082_o_0;
 wire n_13083_o_0;
 wire n_13084_o_0;
 wire n_13085_o_0;
 wire n_13086_o_0;
 wire n_13087_o_0;
 wire n_13088_o_0;
 wire n_13089_o_0;
 wire n_13090_o_0;
 wire n_13091_o_0;
 wire n_13092_o_0;
 wire n_13093_o_0;
 wire n_13094_o_0;
 wire n_13095_o_0;
 wire n_13096_o_0;
 wire n_13097_o_0;
 wire n_13098_o_0;
 wire n_13099_o_0;
 wire n_13100_o_0;
 wire n_13101_o_0;
 wire n_13102_o_0;
 wire n_13103_o_0;

 INVxp67_ASAP7_75t_R clone1 (.A(_00858_),
    .Y(net1));
 INVxp33_ASAP7_75t_R clone10 (.A(n_5489_o_0),
    .Y(net10));
 OAI31xp33_ASAP7_75t_R clone100 (.A1(n_2452_o_0),
    .A2(ld),
    .A3(n_2457_o_0),
    .B(n_2458_o_0),
    .Y(net100));
 A2O1A1Ixp33_ASAP7_75t_R clone101 (.A1(n_2491_o_0),
    .A2(n_2488_o_0),
    .B(ld),
    .C(n_2482_o_0),
    .Y(net101));
 OAI31xp33_ASAP7_75t_R clone102 (.A1(n_2435_o_0),
    .A2(n_2433_o_0),
    .A3(ld),
    .B(n_2436_o_0),
    .Y(net102));
 A2O1A1O1Ixp25_ASAP7_75t_R clone11 (.A1(n_3620_o_0),
    .A2(net),
    .B(n_3621_o_0),
    .C(_00919_),
    .D(n_3622_o_0),
    .Y(net11));
 INVxp33_ASAP7_75t_R clone12 (.A(n_10580_o_0),
    .Y(net12));
 INVxp33_ASAP7_75t_R clone13 (.A(n_1398_o_0),
    .Y(net13));
 INVxp33_ASAP7_75t_R clone14 (.A(n_829_o_0),
    .Y(net14));
 INVxp33_ASAP7_75t_R clone15 (.A(n_829_o_0),
    .Y(net15));
 A2O1A1O1Ixp25_ASAP7_75t_R clone16 (.A1(n_824_o_0),
    .A2(n_825_o_0),
    .B(n_826_o_0),
    .C(n_827_o_0),
    .D(n_828_o_0),
    .Y(net16));
 INVxp33_ASAP7_75t_R clone17 (.A(n_1890_o_0),
    .Y(net17));
 INVxp33_ASAP7_75t_R clone18 (.A(n_1890_o_0),
    .Y(net18));
 A2O1A1Ixp33_ASAP7_75t_R clone19 (.A1(n_8896_o_0),
    .A2(n_8897_o_0),
    .B(n_8898_o_0),
    .C(n_8903_o_0),
    .Y(net19));
 INVx1_ASAP7_75t_R clone2 (.A(_00858_),
    .Y(net2));
 INVxp33_ASAP7_75t_R clone20 (.A(n_1398_o_0),
    .Y(net20));
 A2O1A1O1Ixp25_ASAP7_75t_R clone21 (.A1(_00982_),
    .A2(n_2476_o_0),
    .B(n_2481_o_0),
    .C(n_827_o_0),
    .D(n_2483_o_0),
    .Y(net21));
 NOR2xp33_ASAP7_75t_R clone22 (.A(n_9482_o_0),
    .B(n_9451_o_0),
    .Y(net22));
 NOR2xp33_ASAP7_75t_R clone23 (.A(n_7200_o_0),
    .B(n_7179_o_0),
    .Y(net23));
 A2O1A1O1Ixp25_ASAP7_75t_R clone24 (.A1(net5),
    .A2(_00618_),
    .B(n_10010_o_0),
    .C(_00860_),
    .D(n_10011_o_0),
    .Y(net24));
 A2O1A1O1Ixp25_ASAP7_75t_R clone25 (.A1(net39),
    .A2(n_3670_o_0),
    .B(n_3671_o_0),
    .C(n_2421_o_0),
    .D(n_3672_o_0),
    .Y(net25));
 A2O1A1Ixp33_ASAP7_75t_R clone26 (.A1(n_9473_o_0),
    .A2(n_9474_o_0),
    .B(n_9475_o_0),
    .C(n_9481_o_0),
    .Y(net26));
 O2A1O1Ixp33_ASAP7_75t_R clone27 (.A1(n_3021_o_0),
    .A2(n_4260_o_0),
    .B(n_4316_o_0),
    .C(n_4253_o_0),
    .Y(net27));
 INVxp33_ASAP7_75t_R clone28 (.A(n_1372_o_0),
    .Y(net28));
 A2O1A1Ixp33_ASAP7_75t_R clone29 (.A1(net3),
    .A2(_00492_),
    .B(n_3040_o_0),
    .C(n_3044_o_0),
    .Y(net29));
 INVx1_ASAP7_75t_R clone3 (.A(_00858_),
    .Y(net3));
 O2A1O1Ixp33_ASAP7_75t_R clone30 (.A1(n_3021_o_0),
    .A2(n_3650_o_0),
    .B(n_3652_o_0),
    .C(n_3658_o_0),
    .Y(net30));
 A2O1A1O1Ixp25_ASAP7_75t_R clone31 (.A1(n_1876_o_0),
    .A2(n_1877_o_0),
    .B(n_1878_o_0),
    .C(n_827_o_0),
    .D(n_1879_o_0),
    .Y(net31));
 O2A1O1Ixp33_ASAP7_75t_R clone32 (.A1(n_827_o_0),
    .A2(key[18]),
    .B(n_834_o_0),
    .C(n_835_o_0),
    .Y(net32));
 OAI31xp33_ASAP7_75t_R clone33 (.A1(n_1925_o_0),
    .A2(n_1923_o_0),
    .A3(ld),
    .B(n_1926_o_0),
    .Y(net33));
 A2O1A1Ixp33_ASAP7_75t_R clone34 (.A1(n_7789_o_0),
    .A2(n_7790_o_0),
    .B(n_7777_o_0),
    .C(n_7791_o_0),
    .Y(net34));
 O2A1O1Ixp33_ASAP7_75t_R clone35 (.A1(n_3021_o_0),
    .A2(n_11130_o_0),
    .B(n_11132_o_0),
    .C(n_11135_o_0),
    .Y(net35));
 O2A1O1Ixp33_ASAP7_75t_R clone36 (.A1(n_3097_o_0),
    .A2(net39),
    .B(n_3100_o_0),
    .C(n_3102_o_0),
    .Y(net36));
 A2O1A1Ixp33_ASAP7_75t_R clone37 (.A1(n_11121_o_0),
    .A2(net39),
    .B(n_11123_o_0),
    .C(n_11126_o_0),
    .Y(net37));
 A2O1A1Ixp33_ASAP7_75t_R clone38 (.A1(n_8368_o_0),
    .A2(n_8369_o_0),
    .B(n_8361_o_0),
    .C(n_8362_o_0),
    .Y(net38));
 INVxp33_ASAP7_75t_R clone4 (.A(n_1927_o_0),
    .Y(net4));
 O2A1O1Ixp33_ASAP7_75t_R clone40 (.A1(n_3021_o_0),
    .A2(n_3091_o_0),
    .B(n_3092_o_0),
    .C(n_3076_o_0),
    .Y(net40));
 A2O1A1O1Ixp25_ASAP7_75t_R clone41 (.A1(net39),
    .A2(n_3620_o_0),
    .B(n_3621_o_0),
    .C(n_2399_o_0),
    .D(n_3625_o_0),
    .Y(net41));
 A2O1A1O1Ixp25_ASAP7_75t_R clone42 (.A1(n_824_o_0),
    .A2(n_825_o_0),
    .B(n_826_o_0),
    .C(n_827_o_0),
    .D(n_828_o_0),
    .Y(net42));
 AOI21xp33_ASAP7_75t_R clone43 (.A1(n_10568_o_0),
    .A2(n_10576_o_0),
    .B(n_10579_o_0),
    .Y(net43));
 INVxp33_ASAP7_75t_R clone44 (.A(n_1398_o_0),
    .Y(net44));
 A2O1A1O1Ixp25_ASAP7_75t_R clone45 (.A1(net5),
    .A2(_00581_),
    .B(n_8338_o_0),
    .C(_00901_),
    .D(n_8344_o_0),
    .Y(net45));
 AOI21xp5_ASAP7_75t_R clone46 (.A1(n_7192_o_0),
    .A2(n_7191_o_0),
    .B(n_7195_o_0),
    .Y(net46));
 O2A1O1Ixp33_ASAP7_75t_R clone47 (.A1(n_4192_o_0),
    .A2(net39),
    .B(n_4198_o_0),
    .C(n_4243_o_0),
    .Y(net47));
 A2O1A1Ixp33_ASAP7_75t_R clone48 (.A1(n_8896_o_0),
    .A2(n_8897_o_0),
    .B(n_8898_o_0),
    .C(n_8903_o_0),
    .Y(net48));
 INVx1_ASAP7_75t_R clone5 (.A(_00858_),
    .Y(net5));
 A2O1A1O1Ixp25_ASAP7_75t_R clone50 (.A1(net39),
    .A2(n_3670_o_0),
    .B(n_3671_o_0),
    .C(n_2421_o_0),
    .D(n_3672_o_0),
    .Y(net50));
 A2O1A1O1Ixp25_ASAP7_75t_R clone51 (.A1(net9),
    .A2(_00712_),
    .B(n_4964_o_0),
    .C(_00984_),
    .D(n_4984_o_0),
    .Y(net51));
 OAI31xp33_ASAP7_75t_R clone52 (.A1(ld),
    .A2(n_2410_o_0),
    .A3(n_2413_o_0),
    .B(n_2414_o_0),
    .Y(net52));
 A2O1A1Ixp33_ASAP7_75t_R clone53 (.A1(n_9473_o_0),
    .A2(n_9474_o_0),
    .B(n_9475_o_0),
    .C(n_9481_o_0),
    .Y(net53));
 AOI21xp33_ASAP7_75t_R clone54 (.A1(n_5468_o_0),
    .A2(n_5488_o_0),
    .B(n_5469_o_0),
    .Y(net54));
 AOI21xp33_ASAP7_75t_R clone55 (.A1(n_6604_o_0),
    .A2(n_6610_o_0),
    .B(n_6613_o_0),
    .Y(net55));
 AOI21xp5_ASAP7_75t_R clone56 (.A1(n_10026_o_0),
    .A2(n_10033_o_0),
    .B(n_10036_o_0),
    .Y(net56));
 A2O1A1Ixp33_ASAP7_75t_R clone57 (.A1(n_4918_o_0),
    .A2(net39),
    .B(n_4919_o_0),
    .C(n_4933_o_0),
    .Y(net57));
 O2A1O1Ixp33_ASAP7_75t_R clone58 (.A1(net5),
    .A2(n_11121_o_0),
    .B(n_11125_o_0),
    .C(n_11138_o_0),
    .Y(net58));
 O2A1O1Ixp33_ASAP7_75t_R clone59 (.A1(n_3021_o_0),
    .A2(n_4217_o_0),
    .B(n_4218_o_0),
    .C(n_4225_o_0),
    .Y(net59));
 INVxp33_ASAP7_75t_R clone6 (.A(n_10580_o_0),
    .Y(net6));
 O2A1O1Ixp33_ASAP7_75t_R clone60 (.A1(n_4874_o_0),
    .A2(net39),
    .B(n_4951_o_0),
    .C(n_4872_o_0),
    .Y(net60));
 OAI31xp33_ASAP7_75t_R clone61 (.A1(_00860_),
    .A2(n_10038_o_0),
    .A3(n_10010_o_0),
    .B(n_10039_o_0),
    .Y(net61));
 A2O1A1Ixp33_ASAP7_75t_R clone62 (.A1(n_4190_o_0),
    .A2(net),
    .B(n_4191_o_0),
    .C(n_4199_o_0),
    .Y(net62));
 A2O1A1O1Ixp25_ASAP7_75t_R clone63 (.A1(n_3620_o_0),
    .A2(net39),
    .B(n_3621_o_0),
    .C(_00919_),
    .D(n_3622_o_0),
    .Y(net63));
 A2O1A1O1Ixp25_ASAP7_75t_R clone64 (.A1(n_8885_o_0),
    .A2(net),
    .B(n_8886_o_0),
    .C(_00936_),
    .D(n_8971_o_0),
    .Y(net64));
 AOI21xp5_ASAP7_75t_R clone65 (.A1(n_11146_o_0),
    .A2(n_11140_o_0),
    .B(n_11151_o_0),
    .Y(net65));
 A2O1A1Ixp33_ASAP7_75t_R clone66 (.A1(n_8368_o_0),
    .A2(n_8369_o_0),
    .B(n_8361_o_0),
    .C(n_8362_o_0),
    .Y(net66));
 AOI21xp33_ASAP7_75t_R clone67 (.A1(_00900_),
    .A2(n_8327_o_0),
    .B(n_8331_o_0),
    .Y(net67));
 A2O1A1Ixp33_ASAP7_75t_R clone68 (.A1(n_11121_o_0),
    .A2(net39),
    .B(n_11123_o_0),
    .C(n_11126_o_0),
    .Y(net68));
 O2A1O1Ixp33_ASAP7_75t_R clone69 (.A1(n_4920_o_0),
    .A2(net),
    .B(n_4973_o_0),
    .C(n_4974_o_0),
    .Y(net69));
 INVxp33_ASAP7_75t_R clone7 (.A(n_5489_o_0),
    .Y(net7));
 INVxp33_ASAP7_75t_R clone70 (.A(n_1398_o_0),
    .Y(net70));
 AOI21xp33_ASAP7_75t_R clone71 (.A1(n_827_o_0),
    .A2(n_1396_o_0),
    .B(n_1397_o_0),
    .Y(net71));
 O2A1O1Ixp33_ASAP7_75t_R clone72 (.A1(n_3628_o_0),
    .A2(net),
    .B(n_3636_o_0),
    .C(n_3682_o_0),
    .Y(net72));
 AOI21xp33_ASAP7_75t_R clone73 (.A1(n_8313_o_0),
    .A2(n_8305_o_0),
    .B(n_8317_o_0),
    .Y(net73));
 O2A1O1Ixp33_ASAP7_75t_R clone74 (.A1(n_3021_o_0),
    .A2(n_3650_o_0),
    .B(n_3652_o_0),
    .C(n_3658_o_0),
    .Y(net74));
 A2O1A1O1Ixp25_ASAP7_75t_R clone75 (.A1(_00982_),
    .A2(n_2476_o_0),
    .B(n_2481_o_0),
    .C(n_827_o_0),
    .D(n_2483_o_0),
    .Y(net75));
 A2O1A1O1Ixp25_ASAP7_75t_R clone76 (.A1(net9),
    .A2(_00410_),
    .B(n_11746_o_0),
    .C(_00957_),
    .D(n_11747_o_0),
    .Y(net76));
 A2O1A1O1Ixp25_ASAP7_75t_R clone78 (.A1(_00876_),
    .A2(n_5478_o_0),
    .B(n_5482_o_0),
    .C(n_5459_o_0),
    .D(n_5580_o_0),
    .Y(net78));
 AOI21xp33_ASAP7_75t_R clone79 (.A1(_00973_),
    .A2(n_7165_o_0),
    .B(n_7181_o_0),
    .Y(net79));
 INVxp33_ASAP7_75t_R clone8 (.A(n_1927_o_0),
    .Y(net8));
 A2O1A1Ixp33_ASAP7_75t_R clone82 (.A1(net),
    .A2(n_4217_o_0),
    .B(n_4224_o_0),
    .C(n_4281_o_0),
    .Y(net82));
 AOI21xp33_ASAP7_75t_R clone85 (.A1(n_9519_o_0),
    .A2(n_9511_o_0),
    .B(n_9435_o_0),
    .Y(net85));
 A2O1A1O1Ixp25_ASAP7_75t_R clone86 (.A1(net39),
    .A2(n_3670_o_0),
    .B(n_3671_o_0),
    .C(n_2421_o_0),
    .D(n_3672_o_0),
    .Y(net86));
 A2O1A1Ixp33_ASAP7_75t_R clone89 (.A1(_00964_),
    .A2(n_9444_o_0),
    .B(n_9450_o_0),
    .C(n_9482_o_0),
    .Y(net89));
 INVxp67_ASAP7_75t_R clone9 (.A(_00858_),
    .Y(net9));
 A2O1A1O1Ixp25_ASAP7_75t_R clone90 (.A1(net39),
    .A2(n_3620_o_0),
    .B(n_3621_o_0),
    .C(n_2399_o_0),
    .D(n_3625_o_0),
    .Y(net90));
 A2O1A1O1Ixp25_ASAP7_75t_R clone93 (.A1(n_3620_o_0),
    .A2(net39),
    .B(n_3621_o_0),
    .C(_00919_),
    .D(n_3622_o_0),
    .Y(net93));
 A2O1A1O1Ixp25_ASAP7_75t_R clone94 (.A1(n_3620_o_0),
    .A2(net),
    .B(n_3621_o_0),
    .C(_00919_),
    .D(n_3622_o_0),
    .Y(net94));
 OAI21xp33_ASAP7_75t_R clone95 (.A1(n_4848_o_0),
    .A2(n_2411_o_0),
    .B(n_4953_o_0),
    .Y(net95));
 A2O1A1O1Ixp25_ASAP7_75t_R clone96 (.A1(net9),
    .A2(_00569_),
    .B(n_7775_o_0),
    .C(_00869_),
    .D(n_7778_o_0),
    .Y(net96));
 A2O1A1Ixp33_ASAP7_75t_R clone97 (.A1(n_7789_o_0),
    .A2(n_7790_o_0),
    .B(n_7777_o_0),
    .C(n_7791_o_0),
    .Y(net97));
 INVxp33_ASAP7_75t_R clone98 (.A(n_1890_o_0),
    .Y(net98));
 NAND2xp33_ASAP7_75t_R clone99 (.A(n_1371_o_0),
    .B(n_1368_o_0),
    .Y(net99));
 DFFHQNx1_ASAP7_75t_R \dcnt[0]$_SDFFE_PN0P_  (.CLK(clk),
    .D(n_12874_o_0),
    .QN(_00648_));
 DFFHQNx1_ASAP7_75t_R \dcnt[1]$_SDFFE_PN0P_  (.CLK(clk),
    .D(n_12877_o_0),
    .QN(_00647_));
 DFFHQNx1_ASAP7_75t_R \dcnt[2]$_SDFFE_PP0P_  (.CLK(clk),
    .D(n_12881_o_0),
    .QN(_00645_));
 DFFHQNx1_ASAP7_75t_R \dcnt[3]$_SDFFE_PN0P_  (.CLK(clk),
    .D(n_12879_o_0),
    .QN(_00729_));
 DFFHQNx1_ASAP7_75t_R \done$_DFF_P_  (.CLK(clk),
    .D(n_12241_o_0),
    .QN(_00646_));
 DFFHQNx3_ASAP7_75t_R \ld_r$_DFF_P_  (.CLK(clk),
    .D(ld),
    .QN(_00858_));
 NAND2xp33_ASAP7_75t_R n_1000 (.A(n_877_o_0),
    .B(n_866_o_0),
    .Y(n_1000_o_0));
 XOR2xp5_ASAP7_75t_R n_10000 (.A(_01000_),
    .B(_01001_),
    .Y(n_10000_o_0));
 NOR2xp33_ASAP7_75t_R n_10001 (.A(n_10000_o_0),
    .B(n_9999_o_0),
    .Y(n_10001_o_0));
 NOR2xp33_ASAP7_75t_R n_10002 (.A(_00666_),
    .B(net),
    .Y(n_10002_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10003 (.A1(n_9999_o_0),
    .A2(n_10000_o_0),
    .B(n_10001_o_0),
    .C(net),
    .D(n_10002_o_0),
    .Y(n_10003_o_0));
 XNOR2xp5_ASAP7_75t_R n_10004 (.A(_00865_),
    .B(n_10003_o_0),
    .Y(n_10004_o_0));
 INVx1_ASAP7_75t_R n_10005 (.A(n_10004_o_0),
    .Y(n_10005_o_0));
 NAND2xp33_ASAP7_75t_R n_10006 (.A(n_3046_o_0),
    .B(n_3060_o_0),
    .Y(n_10006_o_0));
 OAI211xp5_ASAP7_75t_R n_10007 (.A1(n_3046_o_0),
    .A2(n_3060_o_0),
    .B(n_10006_o_0),
    .C(n_7697_o_0),
    .Y(n_10007_o_0));
 NOR2xp33_ASAP7_75t_R n_10008 (.A(n_3046_o_0),
    .B(n_3060_o_0),
    .Y(n_10008_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10009 (.A1(n_3046_o_0),
    .A2(n_3060_o_0),
    .B(n_10008_o_0),
    .C(_00642_),
    .Y(n_10009_o_0));
 NAND3xp33_ASAP7_75t_R n_1001 (.A(n_860_o_0),
    .B(n_881_o_0),
    .C(n_878_o_0),
    .Y(n_1001_o_0));
 AOI21xp33_ASAP7_75t_R n_10010 (.A1(n_10007_o_0),
    .A2(n_10009_o_0),
    .B(n_3021_o_0),
    .Y(n_10010_o_0));
 AOI211xp5_ASAP7_75t_R n_10011 (.A1(net1),
    .A2(_00618_),
    .B(n_10010_o_0),
    .C(_00860_),
    .Y(n_10011_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10012 (.A1(net5),
    .A2(_00618_),
    .B(n_10010_o_0),
    .C(_00860_),
    .D(n_10011_o_0),
    .Y(n_10012_o_0));
 NAND2xp33_ASAP7_75t_R n_10013 (.A(n_7762_o_0),
    .B(n_3036_o_0),
    .Y(n_10013_o_0));
 NAND2xp33_ASAP7_75t_R n_10014 (.A(n_3035_o_0),
    .B(n_7759_o_0),
    .Y(n_10014_o_0));
 XNOR2xp5_ASAP7_75t_R n_10015 (.A(_01077_),
    .B(n_3060_o_0),
    .Y(n_10015_o_0));
 AO21x1_ASAP7_75t_R n_10016 (.A1(n_10013_o_0),
    .A2(n_10014_o_0),
    .B(n_10015_o_0),
    .Y(n_10016_o_0));
 XNOR2xp5_ASAP7_75t_R n_10017 (.A(n_3035_o_0),
    .B(n_7762_o_0),
    .Y(n_10017_o_0));
 AOI21xp33_ASAP7_75t_R n_10018 (.A1(n_10015_o_0),
    .A2(n_10017_o_0),
    .B(n_3021_o_0),
    .Y(n_10018_o_0));
 AOI221xp5_ASAP7_75t_R n_10019 (.A1(net9),
    .A2(_00617_),
    .B1(n_10016_o_0),
    .B2(n_10018_o_0),
    .C(_00861_),
    .Y(n_10019_o_0));
 NAND3xp33_ASAP7_75t_R n_1002 (.A(n_935_o_0),
    .B(n_877_o_0),
    .C(n_881_o_0),
    .Y(n_1002_o_0));
 INVx1_ASAP7_75t_R n_10020 (.A(_00617_),
    .Y(n_10020_o_0));
 OAI21xp33_ASAP7_75t_R n_10021 (.A1(n_10017_o_0),
    .A2(n_10015_o_0),
    .B(n_10018_o_0),
    .Y(n_10021_o_0));
 INVx1_ASAP7_75t_R n_10022 (.A(_00861_),
    .Y(n_10022_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10023 (.A1(n_10020_o_0),
    .A2(net),
    .B(n_10021_o_0),
    .C(n_10022_o_0),
    .Y(n_10023_o_0));
 NOR2xp67_ASAP7_75t_R n_10024 (.A(n_10019_o_0),
    .B(n_10023_o_0),
    .Y(n_10024_o_0));
 NOR2xp33_ASAP7_75t_R n_10025 (.A(n_10012_o_0),
    .B(n_10024_o_0),
    .Y(n_10025_o_0));
 INVx1_ASAP7_75t_R n_10026 (.A(_00862_),
    .Y(n_10026_o_0));
 XOR2xp5_ASAP7_75t_R n_10027 (.A(_01078_),
    .B(_01116_),
    .Y(n_10027_o_0));
 NAND2xp33_ASAP7_75t_R n_10028 (.A(_00997_),
    .B(n_10027_o_0),
    .Y(n_10028_o_0));
 OAI21xp33_ASAP7_75t_R n_10029 (.A1(_00997_),
    .A2(n_10027_o_0),
    .B(n_10028_o_0),
    .Y(n_10029_o_0));
 NAND4xp25_ASAP7_75t_R n_1003 (.A(n_1000_o_0),
    .B(n_1001_o_0),
    .C(n_1002_o_0),
    .D(net16),
    .Y(n_1003_o_0));
 OAI211xp5_ASAP7_75t_R n_10030 (.A1(_00997_),
    .A2(n_10027_o_0),
    .B(n_10028_o_0),
    .C(n_7745_o_0),
    .Y(n_10030_o_0));
 INVx1_ASAP7_75t_R n_10031 (.A(n_10030_o_0),
    .Y(n_10031_o_0));
 NOR2xp33_ASAP7_75t_R n_10032 (.A(_00620_),
    .B(net39),
    .Y(n_10032_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10033 (.A1(n_7742_o_0),
    .A2(n_10029_o_0),
    .B(n_10031_o_0),
    .C(net39),
    .D(n_10032_o_0),
    .Y(n_10033_o_0));
 NAND2xp33_ASAP7_75t_R n_10034 (.A(n_7742_o_0),
    .B(n_10029_o_0),
    .Y(n_10034_o_0));
 INVx1_ASAP7_75t_R n_10035 (.A(n_10032_o_0),
    .Y(n_10035_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10036 (.A1(n_10030_o_0),
    .A2(n_10034_o_0),
    .B(n_3021_o_0),
    .C(n_10035_o_0),
    .D(n_10026_o_0),
    .Y(n_10036_o_0));
 AO21x1_ASAP7_75t_R n_10037 (.A1(n_10026_o_0),
    .A2(n_10033_o_0),
    .B(n_10036_o_0),
    .Y(n_10037_o_0));
 AND2x2_ASAP7_75t_R n_10038 (.A(n_3021_o_0),
    .B(_00618_),
    .Y(n_10038_o_0));
 OAI21xp33_ASAP7_75t_R n_10039 (.A1(n_10038_o_0),
    .A2(n_10010_o_0),
    .B(_00860_),
    .Y(n_10039_o_0));
 OAI21xp33_ASAP7_75t_R n_1004 (.A1(n_836_o_0),
    .A2(n_935_o_0),
    .B(n_878_o_0),
    .Y(n_1004_o_0));
 OAI31xp67_ASAP7_75t_R n_10040 (.A1(_00860_),
    .A2(n_10038_o_0),
    .A3(n_10010_o_0),
    .B(n_10039_o_0),
    .Y(n_10040_o_0));
 AOI22xp33_ASAP7_75t_R n_10041 (.A1(n_10018_o_0),
    .A2(n_10016_o_0),
    .B1(n_3021_o_0),
    .B2(_00617_),
    .Y(n_10041_o_0));
 OAI211xp5_ASAP7_75t_R n_10042 (.A1(n_10020_o_0),
    .A2(net39),
    .B(n_10021_o_0),
    .C(n_10022_o_0),
    .Y(n_10042_o_0));
 OAI21x1_ASAP7_75t_R n_10043 (.A1(n_10041_o_0),
    .A2(n_10022_o_0),
    .B(n_10042_o_0),
    .Y(n_10043_o_0));
 AOI21xp33_ASAP7_75t_R n_10044 (.A1(n_10040_o_0),
    .A2(n_10043_o_0),
    .B(n_10037_o_0),
    .Y(n_10044_o_0));
 INVx1_ASAP7_75t_R n_10045 (.A(_00863_),
    .Y(n_10045_o_0));
 XNOR2xp5_ASAP7_75t_R n_10046 (.A(_01079_),
    .B(n_3022_o_0),
    .Y(n_10046_o_0));
 NAND2xp33_ASAP7_75t_R n_10047 (.A(n_10046_o_0),
    .B(n_7727_o_0),
    .Y(n_10047_o_0));
 OAI21xp33_ASAP7_75t_R n_10048 (.A1(n_7727_o_0),
    .A2(n_10046_o_0),
    .B(n_10047_o_0),
    .Y(n_10048_o_0));
 NOR2xp33_ASAP7_75t_R n_10049 (.A(_00668_),
    .B(net77),
    .Y(n_10049_o_0));
 OAI21xp33_ASAP7_75t_R n_1005 (.A1(n_847_o_0),
    .A2(n_864_o_0),
    .B(n_836_o_0),
    .Y(n_1005_o_0));
 AOI21xp33_ASAP7_75t_R n_10050 (.A1(net77),
    .A2(n_10048_o_0),
    .B(n_10049_o_0),
    .Y(n_10050_o_0));
 INVx1_ASAP7_75t_R n_10051 (.A(_01079_),
    .Y(n_10051_o_0));
 NOR2xp33_ASAP7_75t_R n_10052 (.A(n_10051_o_0),
    .B(n_3022_o_0),
    .Y(n_10052_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10053 (.A1(n_3022_o_0),
    .A2(n_10051_o_0),
    .B(n_10052_o_0),
    .C(n_7735_o_0),
    .Y(n_10053_o_0));
 INVx1_ASAP7_75t_R n_10054 (.A(n_10049_o_0),
    .Y(n_10054_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10055 (.A1(n_10053_o_0),
    .A2(n_10047_o_0),
    .B(net3),
    .C(n_10054_o_0),
    .D(n_10045_o_0),
    .Y(n_10055_o_0));
 AOI21x1_ASAP7_75t_R n_10056 (.A1(n_10045_o_0),
    .A2(n_10050_o_0),
    .B(n_10055_o_0),
    .Y(n_10056_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10057 (.A1(n_10025_o_0),
    .A2(n_10037_o_0),
    .B(n_10044_o_0),
    .C(n_10056_o_0),
    .Y(n_10057_o_0));
 AOI21x1_ASAP7_75t_R n_10058 (.A1(n_10026_o_0),
    .A2(n_10033_o_0),
    .B(n_10036_o_0),
    .Y(n_10058_o_0));
 NOR2xp67_ASAP7_75t_R n_10059 (.A(n_10012_o_0),
    .B(n_10043_o_0),
    .Y(n_10059_o_0));
 INVx1_ASAP7_75t_R n_1006 (.A(n_1005_o_0),
    .Y(n_1006_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10060 (.A1(n_10053_o_0),
    .A2(n_10047_o_0),
    .B(net9),
    .C(n_10054_o_0),
    .D(_00863_),
    .Y(n_10060_o_0));
 AOI21xp5_ASAP7_75t_R n_10061 (.A1(_00863_),
    .A2(n_10050_o_0),
    .B(n_10060_o_0),
    .Y(n_10061_o_0));
 OAI21xp33_ASAP7_75t_R n_10062 (.A1(net56),
    .A2(n_10059_o_0),
    .B(n_10061_o_0),
    .Y(n_10062_o_0));
 XNOR2xp5_ASAP7_75t_R n_10063 (.A(_01080_),
    .B(n_3115_o_0),
    .Y(n_10063_o_0));
 XOR2xp5_ASAP7_75t_R n_10064 (.A(n_10063_o_0),
    .B(n_7717_o_0),
    .Y(n_10064_o_0));
 NOR2xp33_ASAP7_75t_R n_10065 (.A(_00667_),
    .B(net39),
    .Y(n_10065_o_0));
 AOI21xp33_ASAP7_75t_R n_10066 (.A1(net),
    .A2(n_10064_o_0),
    .B(n_10065_o_0),
    .Y(n_10066_o_0));
 XNOR2xp5_ASAP7_75t_R n_10067 (.A(_00864_),
    .B(n_10066_o_0),
    .Y(n_10067_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10068 (.A1(n_10022_o_0),
    .A2(n_10041_o_0),
    .B(n_10042_o_0),
    .C(n_10040_o_0),
    .Y(n_10068_o_0));
 NAND2xp33_ASAP7_75t_R n_10069 (.A(n_10058_o_0),
    .B(n_10068_o_0),
    .Y(n_10069_o_0));
 OAI21xp33_ASAP7_75t_R n_1007 (.A1(n_1004_o_0),
    .A2(n_1006_o_0),
    .B(n_960_o_0),
    .Y(n_1007_o_0));
 INVx1_ASAP7_75t_R n_10070 (.A(n_10069_o_0),
    .Y(n_10070_o_0));
 AOI21xp33_ASAP7_75t_R n_10071 (.A1(n_10040_o_0),
    .A2(n_10037_o_0),
    .B(n_10056_o_0),
    .Y(n_10071_o_0));
 INVx1_ASAP7_75t_R n_10072 (.A(n_10071_o_0),
    .Y(n_10072_o_0));
 NAND2xp33_ASAP7_75t_R n_10073 (.A(n_10037_o_0),
    .B(n_10024_o_0),
    .Y(n_10073_o_0));
 OA21x2_ASAP7_75t_R n_10074 (.A1(n_10010_o_0),
    .A2(n_10038_o_0),
    .B(_00860_),
    .Y(n_10074_o_0));
 OAI22xp33_ASAP7_75t_R n_10075 (.A1(n_10019_o_0),
    .A2(n_10023_o_0),
    .B1(n_10074_o_0),
    .B2(n_10011_o_0),
    .Y(n_10075_o_0));
 OAI211xp5_ASAP7_75t_R n_10076 (.A1(n_10043_o_0),
    .A2(n_10040_o_0),
    .B(n_10075_o_0),
    .C(n_10058_o_0),
    .Y(n_10076_o_0));
 AO21x1_ASAP7_75t_R n_10077 (.A1(n_10050_o_0),
    .A2(_00863_),
    .B(n_10060_o_0),
    .Y(n_10077_o_0));
 NAND3xp33_ASAP7_75t_R n_10078 (.A(n_10073_o_0),
    .B(n_10076_o_0),
    .C(n_10077_o_0),
    .Y(n_10078_o_0));
 OAI21xp33_ASAP7_75t_R n_10079 (.A1(n_10070_o_0),
    .A2(n_10072_o_0),
    .B(n_10078_o_0),
    .Y(n_10079_o_0));
 AOI31xp33_ASAP7_75t_R n_1008 (.A1(n_1003_o_0),
    .A2(n_1007_o_0),
    .A3(n_904_o_0),
    .B(n_931_o_0),
    .Y(n_1008_o_0));
 NAND2xp33_ASAP7_75t_R n_10080 (.A(n_10067_o_0),
    .B(n_10079_o_0),
    .Y(n_10080_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10081 (.A1(n_10057_o_0),
    .A2(n_10062_o_0),
    .B(n_10067_o_0),
    .C(n_10080_o_0),
    .Y(n_10081_o_0));
 NAND2xp33_ASAP7_75t_R n_10082 (.A(n_10037_o_0),
    .B(n_10068_o_0),
    .Y(n_10082_o_0));
 NOR3xp33_ASAP7_75t_R n_10083 (.A(n_10037_o_0),
    .B(n_10043_o_0),
    .C(n_10012_o_0),
    .Y(n_10083_o_0));
 INVx1_ASAP7_75t_R n_10084 (.A(n_10083_o_0),
    .Y(n_10084_o_0));
 INVx2_ASAP7_75t_R n_10085 (.A(n_10056_o_0),
    .Y(n_10085_o_0));
 AOI21xp33_ASAP7_75t_R n_10086 (.A1(n_10082_o_0),
    .A2(n_10084_o_0),
    .B(n_10085_o_0),
    .Y(n_10086_o_0));
 OAI21xp5_ASAP7_75t_R n_10087 (.A1(n_10040_o_0),
    .A2(n_10043_o_0),
    .B(n_10075_o_0),
    .Y(n_10087_o_0));
 AOI21xp33_ASAP7_75t_R n_10088 (.A1(n_10037_o_0),
    .A2(n_10087_o_0),
    .B(n_10077_o_0),
    .Y(n_10088_o_0));
 INVx1_ASAP7_75t_R n_10089 (.A(n_10059_o_0),
    .Y(n_10089_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1009 (.A1(n_904_o_0),
    .A2(n_999_o_0),
    .B(n_1008_o_0),
    .C(n_971_o_0),
    .Y(n_1009_o_0));
 NAND2xp33_ASAP7_75t_R n_10090 (.A(n_10058_o_0),
    .B(n_10056_o_0),
    .Y(n_10090_o_0));
 AOI21xp33_ASAP7_75t_R n_10091 (.A1(n_10040_o_0),
    .A2(n_10058_o_0),
    .B(n_10056_o_0),
    .Y(n_10091_o_0));
 NAND3xp33_ASAP7_75t_R n_10092 (.A(n_10024_o_0),
    .B(n_10037_o_0),
    .C(n_10012_o_0),
    .Y(n_10092_o_0));
 INVx1_ASAP7_75t_R n_10093 (.A(n_10067_o_0),
    .Y(n_10093_o_0));
 AOI21xp33_ASAP7_75t_R n_10094 (.A1(n_10091_o_0),
    .A2(n_10092_o_0),
    .B(n_10093_o_0),
    .Y(n_10094_o_0));
 OAI21xp33_ASAP7_75t_R n_10095 (.A1(n_10089_o_0),
    .A2(n_10090_o_0),
    .B(n_10094_o_0),
    .Y(n_10095_o_0));
 OAI31xp33_ASAP7_75t_R n_10096 (.A1(n_10067_o_0),
    .A2(n_10086_o_0),
    .A3(n_10088_o_0),
    .B(n_10095_o_0),
    .Y(n_10096_o_0));
 XOR2xp5_ASAP7_75t_R n_10097 (.A(_00643_),
    .B(_01121_),
    .Y(n_10097_o_0));
 XNOR2xp5_ASAP7_75t_R n_10098 (.A(_01002_),
    .B(n_10097_o_0),
    .Y(n_10098_o_0));
 NOR2xp33_ASAP7_75t_R n_10099 (.A(n_3048_o_0),
    .B(n_10098_o_0),
    .Y(n_10099_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1010 (.A1(n_978_o_0),
    .A2(n_988_o_0),
    .B(n_930_o_0),
    .C(n_1009_o_0),
    .Y(n_1010_o_0));
 NOR2xp33_ASAP7_75t_R n_10100 (.A(_00664_),
    .B(net),
    .Y(n_10100_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10101 (.A1(n_3048_o_0),
    .A2(n_10098_o_0),
    .B(n_10099_o_0),
    .C(net),
    .D(n_10100_o_0),
    .Y(n_10101_o_0));
 XNOR2xp5_ASAP7_75t_R n_10102 (.A(_00867_),
    .B(n_10101_o_0),
    .Y(n_10102_o_0));
 INVx1_ASAP7_75t_R n_10103 (.A(n_10102_o_0),
    .Y(n_10103_o_0));
 OAI21xp33_ASAP7_75t_R n_10104 (.A1(n_10005_o_0),
    .A2(n_10096_o_0),
    .B(n_10103_o_0),
    .Y(n_10104_o_0));
 AOI21xp33_ASAP7_75t_R n_10105 (.A1(n_10005_o_0),
    .A2(n_10081_o_0),
    .B(n_10104_o_0),
    .Y(n_10105_o_0));
 OAI211xp5_ASAP7_75t_R n_10106 (.A1(n_10041_o_0),
    .A2(n_10022_o_0),
    .B(n_10012_o_0),
    .C(n_10042_o_0),
    .Y(n_10106_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10107 (.A1(n_10106_o_0),
    .A2(n_10075_o_0),
    .B(n_10058_o_0),
    .C(n_10085_o_0),
    .Y(n_10107_o_0));
 OAI21xp33_ASAP7_75t_R n_10108 (.A1(n_10040_o_0),
    .A2(n_10043_o_0),
    .B(n_10058_o_0),
    .Y(n_10108_o_0));
 INVx1_ASAP7_75t_R n_10109 (.A(n_10108_o_0),
    .Y(n_10109_o_0));
 OAI31xp33_ASAP7_75t_R n_1011 (.A1(n_932_o_0),
    .A2(n_963_o_0),
    .A3(n_972_o_0),
    .B(n_1010_o_0),
    .Y(n_1011_o_0));
 AOI21xp33_ASAP7_75t_R n_10110 (.A1(n_10040_o_0),
    .A2(n_10037_o_0),
    .B(n_10061_o_0),
    .Y(n_10110_o_0));
 NOR2xp33_ASAP7_75t_R n_10111 (.A(n_10012_o_0),
    .B(n_10043_o_0),
    .Y(n_10111_o_0));
 INVx1_ASAP7_75t_R n_10112 (.A(n_10111_o_0),
    .Y(n_10112_o_0));
 INVx1_ASAP7_75t_R n_10113 (.A(_00864_),
    .Y(n_10113_o_0));
 AO21x1_ASAP7_75t_R n_10114 (.A1(n_10064_o_0),
    .A2(net),
    .B(n_10065_o_0),
    .Y(n_10114_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10115 (.A1(n_10064_o_0),
    .A2(net),
    .B(n_10065_o_0),
    .C(n_10113_o_0),
    .Y(n_10115_o_0));
 OAI21xp5_ASAP7_75t_R n_10116 (.A1(n_10113_o_0),
    .A2(n_10114_o_0),
    .B(n_10115_o_0),
    .Y(n_10116_o_0));
 AOI21xp33_ASAP7_75t_R n_10117 (.A1(n_10110_o_0),
    .A2(n_10112_o_0),
    .B(n_10116_o_0),
    .Y(n_10117_o_0));
 NAND3xp33_ASAP7_75t_R n_10118 (.A(n_10024_o_0),
    .B(n_10040_o_0),
    .C(n_10058_o_0),
    .Y(n_10118_o_0));
 OAI21xp33_ASAP7_75t_R n_10119 (.A1(n_10012_o_0),
    .A2(n_10043_o_0),
    .B(n_10037_o_0),
    .Y(n_10119_o_0));
 AOI21xp33_ASAP7_75t_R n_1012 (.A1(n_836_o_0),
    .A2(n_913_o_0),
    .B(n_877_o_0),
    .Y(n_1012_o_0));
 AOI21xp33_ASAP7_75t_R n_10120 (.A1(net61),
    .A2(net56),
    .B(n_10061_o_0),
    .Y(n_10120_o_0));
 AOI31xp33_ASAP7_75t_R n_10121 (.A1(n_10085_o_0),
    .A2(n_10118_o_0),
    .A3(n_10119_o_0),
    .B(n_10120_o_0),
    .Y(n_10121_o_0));
 AO21x1_ASAP7_75t_R n_10122 (.A1(n_10121_o_0),
    .A2(n_10067_o_0),
    .B(n_10004_o_0),
    .Y(n_10122_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10123 (.A1(n_10107_o_0),
    .A2(n_10109_o_0),
    .B(n_10117_o_0),
    .C(n_10122_o_0),
    .Y(n_10123_o_0));
 NAND3xp33_ASAP7_75t_R n_10124 (.A(n_10037_o_0),
    .B(n_10043_o_0),
    .C(n_10040_o_0),
    .Y(n_10124_o_0));
 NAND2xp33_ASAP7_75t_R n_10125 (.A(n_10058_o_0),
    .B(n_10043_o_0),
    .Y(n_10125_o_0));
 AO21x1_ASAP7_75t_R n_10126 (.A1(n_10124_o_0),
    .A2(n_10125_o_0),
    .B(n_10085_o_0),
    .Y(n_10126_o_0));
 NAND2xp33_ASAP7_75t_R n_10127 (.A(n_10040_o_0),
    .B(n_10058_o_0),
    .Y(n_10127_o_0));
 OAI21xp33_ASAP7_75t_R n_10128 (.A1(n_10043_o_0),
    .A2(n_10127_o_0),
    .B(n_10077_o_0),
    .Y(n_10128_o_0));
 NOR2xp33_ASAP7_75t_R n_10129 (.A(n_10058_o_0),
    .B(n_10024_o_0),
    .Y(n_10129_o_0));
 OAI21xp33_ASAP7_75t_R n_1013 (.A1(n_889_o_0),
    .A2(net32),
    .B(n_1012_o_0),
    .Y(n_1013_o_0));
 OAI211xp5_ASAP7_75t_R n_10130 (.A1(n_10024_o_0),
    .A2(net56),
    .B(n_10061_o_0),
    .C(net24),
    .Y(n_10130_o_0));
 OA211x2_ASAP7_75t_R n_10131 (.A1(n_10128_o_0),
    .A2(n_10129_o_0),
    .B(n_10093_o_0),
    .C(n_10130_o_0),
    .Y(n_10131_o_0));
 AOI211xp5_ASAP7_75t_R n_10132 (.A1(n_10094_o_0),
    .A2(n_10126_o_0),
    .B(n_10131_o_0),
    .C(n_10005_o_0),
    .Y(n_10132_o_0));
 NOR3xp33_ASAP7_75t_R n_10133 (.A(n_10123_o_0),
    .B(n_10132_o_0),
    .C(n_10103_o_0),
    .Y(n_10133_o_0));
 NAND2xp33_ASAP7_75t_R n_10134 (.A(n_10012_o_0),
    .B(n_10058_o_0),
    .Y(n_10134_o_0));
 AOI21xp33_ASAP7_75t_R n_10135 (.A1(n_10037_o_0),
    .A2(n_10087_o_0),
    .B(n_10085_o_0),
    .Y(n_10135_o_0));
 OAI21xp33_ASAP7_75t_R n_10136 (.A1(n_10043_o_0),
    .A2(n_10134_o_0),
    .B(n_10135_o_0),
    .Y(n_10136_o_0));
 NAND2xp33_ASAP7_75t_R n_10137 (.A(n_10012_o_0),
    .B(n_10043_o_0),
    .Y(n_10137_o_0));
 AOI21xp33_ASAP7_75t_R n_10138 (.A1(net56),
    .A2(n_10025_o_0),
    .B(n_10056_o_0),
    .Y(n_10138_o_0));
 OAI21xp33_ASAP7_75t_R n_10139 (.A1(n_10137_o_0),
    .A2(net56),
    .B(n_10138_o_0),
    .Y(n_10139_o_0));
 OAI31xp33_ASAP7_75t_R n_1014 (.A1(n_935_o_0),
    .A2(net32),
    .A3(n_878_o_0),
    .B(n_1013_o_0),
    .Y(n_1014_o_0));
 NAND2xp33_ASAP7_75t_R n_10140 (.A(n_10040_o_0),
    .B(n_10043_o_0),
    .Y(n_10140_o_0));
 AOI21xp33_ASAP7_75t_R n_10141 (.A1(n_10037_o_0),
    .A2(n_10012_o_0),
    .B(n_10061_o_0),
    .Y(n_10141_o_0));
 NAND2xp33_ASAP7_75t_R n_10142 (.A(n_10140_o_0),
    .B(n_10141_o_0),
    .Y(n_10142_o_0));
 NAND2xp33_ASAP7_75t_R n_10143 (.A(net24),
    .B(n_10058_o_0),
    .Y(n_10143_o_0));
 OAI211xp5_ASAP7_75t_R n_10144 (.A1(n_10043_o_0),
    .A2(net24),
    .B(n_10085_o_0),
    .C(n_10143_o_0),
    .Y(n_10144_o_0));
 AND2x2_ASAP7_75t_R n_10145 (.A(n_10142_o_0),
    .B(n_10144_o_0),
    .Y(n_10145_o_0));
 INVx1_ASAP7_75t_R n_10146 (.A(n_10116_o_0),
    .Y(n_10146_o_0));
 AOI321xp33_ASAP7_75t_R n_10147 (.A1(n_10136_o_0),
    .A2(n_10139_o_0),
    .A3(n_10067_o_0),
    .B1(n_10145_o_0),
    .B2(n_10146_o_0),
    .C(n_10004_o_0),
    .Y(n_10147_o_0));
 NAND2xp33_ASAP7_75t_R n_10148 (.A(_00865_),
    .B(n_10003_o_0),
    .Y(n_10148_o_0));
 OAI21xp33_ASAP7_75t_R n_10149 (.A1(_00865_),
    .A2(n_10003_o_0),
    .B(n_10148_o_0),
    .Y(n_10149_o_0));
 NOR3xp33_ASAP7_75t_R n_1015 (.A(n_938_o_0),
    .B(n_877_o_0),
    .C(n_952_o_0),
    .Y(n_1015_o_0));
 INVx1_ASAP7_75t_R n_10150 (.A(n_10149_o_0),
    .Y(n_10150_o_0));
 INVx1_ASAP7_75t_R n_10151 (.A(n_10124_o_0),
    .Y(n_10151_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10152 (.A1(n_10041_o_0),
    .A2(n_10022_o_0),
    .B(n_10042_o_0),
    .C(n_10012_o_0),
    .Y(n_10152_o_0));
 AOI211xp5_ASAP7_75t_R n_10153 (.A1(n_10012_o_0),
    .A2(n_10024_o_0),
    .B(n_10152_o_0),
    .C(n_10056_o_0),
    .Y(n_10153_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10154 (.A1(n_10045_o_0),
    .A2(n_10050_o_0),
    .B(n_10055_o_0),
    .C(n_10058_o_0),
    .Y(n_10154_o_0));
 AOI21xp33_ASAP7_75t_R n_10155 (.A1(n_10075_o_0),
    .A2(n_10106_o_0),
    .B(n_10154_o_0),
    .Y(n_10155_o_0));
 NAND2xp33_ASAP7_75t_R n_10156 (.A(n_10040_o_0),
    .B(n_10043_o_0),
    .Y(n_10156_o_0));
 OAI22xp33_ASAP7_75t_R n_10157 (.A1(n_10153_o_0),
    .A2(n_10155_o_0),
    .B1(n_10156_o_0),
    .B2(n_10037_o_0),
    .Y(n_10157_o_0));
 OAI31xp33_ASAP7_75t_R n_10158 (.A1(n_10070_o_0),
    .A2(n_10061_o_0),
    .A3(n_10151_o_0),
    .B(n_10157_o_0),
    .Y(n_10158_o_0));
 NAND3xp33_ASAP7_75t_R n_10159 (.A(n_10106_o_0),
    .B(n_10037_o_0),
    .C(n_10075_o_0),
    .Y(n_10159_o_0));
 AOI31xp33_ASAP7_75t_R n_1016 (.A1(n_877_o_0),
    .A2(n_881_o_0),
    .A3(n_957_o_0),
    .B(n_1015_o_0),
    .Y(n_1016_o_0));
 OAI21xp33_ASAP7_75t_R n_10160 (.A1(n_10043_o_0),
    .A2(n_10037_o_0),
    .B(n_10056_o_0),
    .Y(n_10160_o_0));
 INVx1_ASAP7_75t_R n_10161 (.A(n_10160_o_0),
    .Y(n_10161_o_0));
 AOI21xp33_ASAP7_75t_R n_10162 (.A1(n_10058_o_0),
    .A2(n_10087_o_0),
    .B(n_10077_o_0),
    .Y(n_10162_o_0));
 AOI211xp5_ASAP7_75t_R n_10163 (.A1(n_10159_o_0),
    .A2(n_10161_o_0),
    .B(n_10162_o_0),
    .C(n_10067_o_0),
    .Y(n_10163_o_0));
 AOI21xp33_ASAP7_75t_R n_10164 (.A1(n_10116_o_0),
    .A2(n_10158_o_0),
    .B(n_10163_o_0),
    .Y(n_10164_o_0));
 OAI21xp33_ASAP7_75t_R n_10165 (.A1(n_10150_o_0),
    .A2(n_10164_o_0),
    .B(n_10102_o_0),
    .Y(n_10165_o_0));
 NOR3xp33_ASAP7_75t_R n_10166 (.A(n_10043_o_0),
    .B(n_10058_o_0),
    .C(n_10012_o_0),
    .Y(n_10166_o_0));
 OAI21xp33_ASAP7_75t_R n_10167 (.A1(n_10037_o_0),
    .A2(n_10068_o_0),
    .B(n_10061_o_0),
    .Y(n_10167_o_0));
 NOR2xp33_ASAP7_75t_R n_10168 (.A(n_10166_o_0),
    .B(n_10167_o_0),
    .Y(n_10168_o_0));
 AOI211xp5_ASAP7_75t_R n_10169 (.A1(n_10056_o_0),
    .A2(n_10151_o_0),
    .B(n_10168_o_0),
    .C(n_10146_o_0),
    .Y(n_10169_o_0));
 AOI21xp33_ASAP7_75t_R n_1017 (.A1(n_904_o_0),
    .A2(n_1016_o_0),
    .B(n_891_o_0),
    .Y(n_1017_o_0));
 NAND2xp33_ASAP7_75t_R n_10170 (.A(n_10037_o_0),
    .B(n_10085_o_0),
    .Y(n_10170_o_0));
 AOI31xp33_ASAP7_75t_R n_10171 (.A1(n_10043_o_0),
    .A2(n_10058_o_0),
    .A3(net24),
    .B(n_10061_o_0),
    .Y(n_10171_o_0));
 NAND3xp33_ASAP7_75t_R n_10172 (.A(n_10024_o_0),
    .B(n_10037_o_0),
    .C(n_10040_o_0),
    .Y(n_10172_o_0));
 AOI21xp33_ASAP7_75t_R n_10173 (.A1(n_10171_o_0),
    .A2(n_10172_o_0),
    .B(n_10116_o_0),
    .Y(n_10173_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10174 (.A1(n_10170_o_0),
    .A2(n_10156_o_0),
    .B(n_10173_o_0),
    .C(n_10004_o_0),
    .Y(n_10174_o_0));
 INVx1_ASAP7_75t_R n_10175 (.A(n_10174_o_0),
    .Y(n_10175_o_0));
 INVx1_ASAP7_75t_R n_10176 (.A(n_10091_o_0),
    .Y(n_10176_o_0));
 OAI21xp33_ASAP7_75t_R n_10177 (.A1(n_10012_o_0),
    .A2(n_10043_o_0),
    .B(n_10058_o_0),
    .Y(n_10177_o_0));
 NAND3xp33_ASAP7_75t_R n_10178 (.A(n_10043_o_0),
    .B(n_10040_o_0),
    .C(n_10058_o_0),
    .Y(n_10178_o_0));
 INVx1_ASAP7_75t_R n_10179 (.A(n_10178_o_0),
    .Y(n_10179_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1018 (.A1(n_903_o_0),
    .A2(n_1014_o_0),
    .B(net15),
    .C(n_1017_o_0),
    .Y(n_1018_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10180 (.A1(n_10172_o_0),
    .A2(n_10177_o_0),
    .B(n_10179_o_0),
    .C(n_10077_o_0),
    .D(n_10093_o_0),
    .Y(n_10180_o_0));
 OAI21xp33_ASAP7_75t_R n_10181 (.A1(n_10176_o_0),
    .A2(n_10151_o_0),
    .B(n_10180_o_0),
    .Y(n_10181_o_0));
 NOR2xp33_ASAP7_75t_R n_10182 (.A(n_10058_o_0),
    .B(n_10043_o_0),
    .Y(n_10182_o_0));
 AOI21xp33_ASAP7_75t_R n_10183 (.A1(n_10061_o_0),
    .A2(n_10182_o_0),
    .B(n_10067_o_0),
    .Y(n_10183_o_0));
 OAI21xp33_ASAP7_75t_R n_10184 (.A1(n_10085_o_0),
    .A2(n_10076_o_0),
    .B(n_10183_o_0),
    .Y(n_10184_o_0));
 AOI31xp33_ASAP7_75t_R n_10185 (.A1(n_10004_o_0),
    .A2(n_10181_o_0),
    .A3(n_10184_o_0),
    .B(n_10102_o_0),
    .Y(n_10185_o_0));
 OAI21xp33_ASAP7_75t_R n_10186 (.A1(n_10169_o_0),
    .A2(n_10175_o_0),
    .B(n_10185_o_0),
    .Y(n_10186_o_0));
 NAND2xp33_ASAP7_75t_R n_10187 (.A(_00866_),
    .B(n_9995_o_0),
    .Y(n_10187_o_0));
 OAI21xp33_ASAP7_75t_R n_10188 (.A1(_00866_),
    .A2(n_9995_o_0),
    .B(n_10187_o_0),
    .Y(n_10188_o_0));
 OAI211xp5_ASAP7_75t_R n_10189 (.A1(n_10147_o_0),
    .A2(n_10165_o_0),
    .B(n_10186_o_0),
    .C(n_10188_o_0),
    .Y(n_10189_o_0));
 OAI21xp33_ASAP7_75t_R n_1019 (.A1(n_847_o_0),
    .A2(n_864_o_0),
    .B(n_958_o_0),
    .Y(n_1019_o_0));
 OAI31xp33_ASAP7_75t_R n_10190 (.A1(n_9997_o_0),
    .A2(n_10105_o_0),
    .A3(n_10133_o_0),
    .B(n_10189_o_0),
    .Y(n_10190_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10191 (.A1(n_10037_o_0),
    .A2(n_10156_o_0),
    .B(n_10141_o_0),
    .C(n_10149_o_0),
    .Y(n_10191_o_0));
 AOI211xp5_ASAP7_75t_R n_10192 (.A1(n_10037_o_0),
    .A2(net24),
    .B(n_10043_o_0),
    .C(n_10056_o_0),
    .Y(n_10192_o_0));
 INVx1_ASAP7_75t_R n_10193 (.A(n_10192_o_0),
    .Y(n_10193_o_0));
 INVx1_ASAP7_75t_R n_10194 (.A(n_10092_o_0),
    .Y(n_10194_o_0));
 INVx1_ASAP7_75t_R n_10195 (.A(n_10127_o_0),
    .Y(n_10195_o_0));
 OAI31xp33_ASAP7_75t_R n_10196 (.A1(n_10061_o_0),
    .A2(n_10194_o_0),
    .A3(n_10195_o_0),
    .B(n_10107_o_0),
    .Y(n_10196_o_0));
 OAI21xp33_ASAP7_75t_R n_10197 (.A1(n_10005_o_0),
    .A2(n_10196_o_0),
    .B(n_10116_o_0),
    .Y(n_10197_o_0));
 AOI21xp33_ASAP7_75t_R n_10198 (.A1(n_10191_o_0),
    .A2(n_10193_o_0),
    .B(n_10197_o_0),
    .Y(n_10198_o_0));
 INVx1_ASAP7_75t_R n_10199 (.A(n_10134_o_0),
    .Y(n_10199_o_0));
 OAI21xp33_ASAP7_75t_R n_1020 (.A1(n_991_o_0),
    .A2(n_934_o_0),
    .B(n_1019_o_0),
    .Y(n_1020_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10200 (.A1(n_10106_o_0),
    .A2(n_10075_o_0),
    .B(n_10037_o_0),
    .C(n_10061_o_0),
    .Y(n_10200_o_0));
 OAI21xp33_ASAP7_75t_R n_10201 (.A1(n_10200_o_0),
    .A2(n_10151_o_0),
    .B(n_10150_o_0),
    .Y(n_10201_o_0));
 AOI21xp33_ASAP7_75t_R n_10202 (.A1(n_10199_o_0),
    .A2(n_10077_o_0),
    .B(n_10201_o_0),
    .Y(n_10202_o_0));
 NOR2xp33_ASAP7_75t_R n_10203 (.A(n_10058_o_0),
    .B(n_10061_o_0),
    .Y(n_10203_o_0));
 NAND2xp33_ASAP7_75t_R n_10204 (.A(n_10203_o_0),
    .B(n_10025_o_0),
    .Y(n_10204_o_0));
 INVx1_ASAP7_75t_R n_10205 (.A(n_10087_o_0),
    .Y(n_10205_o_0));
 NOR3xp33_ASAP7_75t_R n_10206 (.A(n_10037_o_0),
    .B(n_10043_o_0),
    .C(n_10040_o_0),
    .Y(n_10206_o_0));
 AOI211xp5_ASAP7_75t_R n_10207 (.A1(n_10205_o_0),
    .A2(n_10037_o_0),
    .B(n_10056_o_0),
    .C(n_10206_o_0),
    .Y(n_10207_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10208 (.A1(n_10024_o_0),
    .A2(net24),
    .B(n_10058_o_0),
    .C(n_10056_o_0),
    .Y(n_10208_o_0));
 AOI21xp33_ASAP7_75t_R n_10209 (.A1(net56),
    .A2(n_10156_o_0),
    .B(n_10208_o_0),
    .Y(n_10209_o_0));
 AOI211xp5_ASAP7_75t_R n_1021 (.A1(n_881_o_0),
    .A2(n_889_o_0),
    .B(n_984_o_0),
    .C(n_877_o_0),
    .Y(n_1021_o_0));
 OAI31xp33_ASAP7_75t_R n_10210 (.A1(n_10005_o_0),
    .A2(n_10207_o_0),
    .A3(n_10209_o_0),
    .B(n_10093_o_0),
    .Y(n_10210_o_0));
 AOI21xp33_ASAP7_75t_R n_10211 (.A1(n_10202_o_0),
    .A2(n_10204_o_0),
    .B(n_10210_o_0),
    .Y(n_10211_o_0));
 NOR3xp33_ASAP7_75t_R n_10212 (.A(n_10198_o_0),
    .B(n_10211_o_0),
    .C(n_10103_o_0),
    .Y(n_10212_o_0));
 AOI21xp33_ASAP7_75t_R n_10213 (.A1(n_10037_o_0),
    .A2(n_10205_o_0),
    .B(n_10206_o_0),
    .Y(n_10213_o_0));
 NAND2xp33_ASAP7_75t_R n_10214 (.A(n_10056_o_0),
    .B(n_10059_o_0),
    .Y(n_10214_o_0));
 INVx1_ASAP7_75t_R n_10215 (.A(n_10214_o_0),
    .Y(n_10215_o_0));
 AOI22xp33_ASAP7_75t_R n_10216 (.A1(n_10213_o_0),
    .A2(n_10085_o_0),
    .B1(n_10037_o_0),
    .B2(n_10215_o_0),
    .Y(n_10216_o_0));
 NOR3xp33_ASAP7_75t_R n_10217 (.A(n_10216_o_0),
    .B(n_10149_o_0),
    .C(n_10146_o_0),
    .Y(n_10217_o_0));
 NOR2xp33_ASAP7_75t_R n_10218 (.A(n_10012_o_0),
    .B(n_10058_o_0),
    .Y(n_10218_o_0));
 NOR2xp33_ASAP7_75t_R n_10219 (.A(n_10040_o_0),
    .B(n_10043_o_0),
    .Y(n_10219_o_0));
 OAI31xp33_ASAP7_75t_R n_1022 (.A1(n_878_o_0),
    .A2(n_861_o_0),
    .A3(n_994_o_0),
    .B(net42),
    .Y(n_1022_o_0));
 OAI21xp33_ASAP7_75t_R n_10220 (.A1(n_10037_o_0),
    .A2(n_10205_o_0),
    .B(n_10141_o_0),
    .Y(n_10220_o_0));
 OAI31xp33_ASAP7_75t_R n_10221 (.A1(n_10056_o_0),
    .A2(n_10218_o_0),
    .A3(n_10219_o_0),
    .B(n_10220_o_0),
    .Y(n_10221_o_0));
 NOR3xp33_ASAP7_75t_R n_10222 (.A(n_10221_o_0),
    .B(n_10150_o_0),
    .C(n_10146_o_0),
    .Y(n_10222_o_0));
 NAND2xp33_ASAP7_75t_R n_10223 (.A(_00867_),
    .B(n_10101_o_0),
    .Y(n_10223_o_0));
 OAI21xp33_ASAP7_75t_R n_10224 (.A1(_00867_),
    .A2(n_10101_o_0),
    .B(n_10223_o_0),
    .Y(n_10224_o_0));
 INVx1_ASAP7_75t_R n_10225 (.A(n_10219_o_0),
    .Y(n_10225_o_0));
 AOI211xp5_ASAP7_75t_R n_10226 (.A1(net56),
    .A2(net61),
    .B(n_10056_o_0),
    .C(n_10043_o_0),
    .Y(n_10226_o_0));
 AOI21xp33_ASAP7_75t_R n_10227 (.A1(n_10203_o_0),
    .A2(n_10225_o_0),
    .B(n_10226_o_0),
    .Y(n_10227_o_0));
 OAI211xp5_ASAP7_75t_R n_10228 (.A1(n_10043_o_0),
    .A2(net56),
    .B(net61),
    .C(n_10056_o_0),
    .Y(n_10228_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10229 (.A1(n_10083_o_0),
    .A2(n_10107_o_0),
    .B(n_10228_o_0),
    .C(n_10005_o_0),
    .Y(n_10229_o_0));
 OAI21xp33_ASAP7_75t_R n_1023 (.A1(n_1021_o_0),
    .A2(n_1022_o_0),
    .B(n_903_o_0),
    .Y(n_1023_o_0));
 AOI211xp5_ASAP7_75t_R n_10230 (.A1(n_10150_o_0),
    .A2(n_10227_o_0),
    .B(n_10229_o_0),
    .C(n_10067_o_0),
    .Y(n_10230_o_0));
 NOR4xp25_ASAP7_75t_R n_10231 (.A(n_10217_o_0),
    .B(n_10222_o_0),
    .C(n_10224_o_0),
    .D(n_10230_o_0),
    .Y(n_10231_o_0));
 NOR2xp33_ASAP7_75t_R n_10232 (.A(n_10037_o_0),
    .B(n_10024_o_0),
    .Y(n_10232_o_0));
 NAND2xp33_ASAP7_75t_R n_10233 (.A(n_10171_o_0),
    .B(n_10092_o_0),
    .Y(n_10233_o_0));
 OAI31xp33_ASAP7_75t_R n_10234 (.A1(n_10056_o_0),
    .A2(n_10150_o_0),
    .A3(n_10232_o_0),
    .B(n_10233_o_0),
    .Y(n_10234_o_0));
 OAI21xp33_ASAP7_75t_R n_10235 (.A1(net61),
    .A2(n_10058_o_0),
    .B(n_10161_o_0),
    .Y(n_10235_o_0));
 NAND3xp33_ASAP7_75t_R n_10236 (.A(n_10235_o_0),
    .B(n_10193_o_0),
    .C(n_10004_o_0),
    .Y(n_10236_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10237 (.A1(n_10037_o_0),
    .A2(n_10156_o_0),
    .B(n_10110_o_0),
    .C(n_10149_o_0),
    .Y(n_10237_o_0));
 NAND3xp33_ASAP7_75t_R n_10238 (.A(n_10092_o_0),
    .B(n_10118_o_0),
    .C(n_10085_o_0),
    .Y(n_10238_o_0));
 AOI21xp33_ASAP7_75t_R n_10239 (.A1(n_10237_o_0),
    .A2(n_10238_o_0),
    .B(n_10067_o_0),
    .Y(n_10239_o_0));
 AOI21xp33_ASAP7_75t_R n_1024 (.A1(net15),
    .A2(n_1020_o_0),
    .B(n_1023_o_0),
    .Y(n_1024_o_0));
 AO21x1_ASAP7_75t_R n_10240 (.A1(n_10236_o_0),
    .A2(n_10239_o_0),
    .B(n_10103_o_0),
    .Y(n_10240_o_0));
 AOI21xp33_ASAP7_75t_R n_10241 (.A1(n_10058_o_0),
    .A2(n_10024_o_0),
    .B(n_10056_o_0),
    .Y(n_10241_o_0));
 NOR2xp33_ASAP7_75t_R n_10242 (.A(n_10058_o_0),
    .B(n_10024_o_0),
    .Y(n_10242_o_0));
 AOI311xp33_ASAP7_75t_R n_10243 (.A1(net56),
    .A2(n_10056_o_0),
    .A3(n_10059_o_0),
    .B(n_10241_o_0),
    .C(n_10242_o_0),
    .Y(n_10243_o_0));
 INVx1_ASAP7_75t_R n_10244 (.A(n_10088_o_0),
    .Y(n_10244_o_0));
 NOR2xp33_ASAP7_75t_R n_10245 (.A(n_10012_o_0),
    .B(n_10037_o_0),
    .Y(n_10245_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10246 (.A1(n_10075_o_0),
    .A2(net61),
    .B(n_10058_o_0),
    .C(n_10056_o_0),
    .Y(n_10246_o_0));
 OAI22xp33_ASAP7_75t_R n_10247 (.A1(n_10244_o_0),
    .A2(n_10245_o_0),
    .B1(n_10246_o_0),
    .B2(n_10199_o_0),
    .Y(n_10247_o_0));
 OAI21xp33_ASAP7_75t_R n_10248 (.A1(n_10004_o_0),
    .A2(n_10247_o_0),
    .B(n_10146_o_0),
    .Y(n_10248_o_0));
 NAND3xp33_ASAP7_75t_R n_10249 (.A(n_10073_o_0),
    .B(n_10140_o_0),
    .C(n_10077_o_0),
    .Y(n_10249_o_0));
 INVx1_ASAP7_75t_R n_1025 (.A(n_941_o_0),
    .Y(n_1025_o_0));
 OAI21xp33_ASAP7_75t_R n_10250 (.A1(n_10111_o_0),
    .A2(n_10154_o_0),
    .B(n_10249_o_0),
    .Y(n_10250_o_0));
 OAI21xp33_ASAP7_75t_R n_10251 (.A1(n_10040_o_0),
    .A2(n_10043_o_0),
    .B(n_10037_o_0),
    .Y(n_10251_o_0));
 AOI21xp33_ASAP7_75t_R n_10252 (.A1(n_10251_o_0),
    .A2(n_10162_o_0),
    .B(n_10150_o_0),
    .Y(n_10252_o_0));
 INVx1_ASAP7_75t_R n_10253 (.A(n_10166_o_0),
    .Y(n_10253_o_0));
 OAI211xp5_ASAP7_75t_R n_10254 (.A1(n_10059_o_0),
    .A2(n_10037_o_0),
    .B(n_10253_o_0),
    .C(n_10056_o_0),
    .Y(n_10254_o_0));
 AOI21xp33_ASAP7_75t_R n_10255 (.A1(n_10252_o_0),
    .A2(n_10254_o_0),
    .B(n_10093_o_0),
    .Y(n_10255_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10256 (.A1(n_10004_o_0),
    .A2(n_10250_o_0),
    .B(n_10255_o_0),
    .C(n_10102_o_0),
    .Y(n_10256_o_0));
 INVx1_ASAP7_75t_R n_10257 (.A(n_9997_o_0),
    .Y(n_10257_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10258 (.A1(n_10149_o_0),
    .A2(n_10243_o_0),
    .B(n_10248_o_0),
    .C(n_10256_o_0),
    .D(n_10257_o_0),
    .Y(n_10258_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10259 (.A1(n_10116_o_0),
    .A2(n_10234_o_0),
    .B(n_10240_o_0),
    .C(n_10258_o_0),
    .Y(n_10259_o_0));
 NAND2xp33_ASAP7_75t_R n_1026 (.A(n_944_o_0),
    .B(n_937_o_0),
    .Y(n_1026_o_0));
 OAI31xp33_ASAP7_75t_R n_10260 (.A1(n_9997_o_0),
    .A2(n_10212_o_0),
    .A3(n_10231_o_0),
    .B(n_10259_o_0),
    .Y(n_10260_o_0));
 INVx1_ASAP7_75t_R n_10261 (.A(n_10125_o_0),
    .Y(n_10261_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10262 (.A1(n_10072_o_0),
    .A2(n_10261_o_0),
    .B(n_10078_o_0),
    .C(n_10004_o_0),
    .Y(n_10262_o_0));
 NOR2xp33_ASAP7_75t_R n_10263 (.A(n_10058_o_0),
    .B(n_10043_o_0),
    .Y(n_10263_o_0));
 NOR2xp33_ASAP7_75t_R n_10264 (.A(n_10044_o_0),
    .B(n_10263_o_0),
    .Y(n_10264_o_0));
 OA211x2_ASAP7_75t_R n_10265 (.A1(n_10068_o_0),
    .A2(net56),
    .B(n_10076_o_0),
    .C(n_10085_o_0),
    .Y(n_10265_o_0));
 AOI211xp5_ASAP7_75t_R n_10266 (.A1(n_10077_o_0),
    .A2(n_10264_o_0),
    .B(n_10265_o_0),
    .C(n_10005_o_0),
    .Y(n_10266_o_0));
 AOI22xp33_ASAP7_75t_R n_10267 (.A1(n_10056_o_0),
    .A2(n_10182_o_0),
    .B1(n_10162_o_0),
    .B2(n_10253_o_0),
    .Y(n_10267_o_0));
 NAND3xp33_ASAP7_75t_R n_10268 (.A(n_10073_o_0),
    .B(n_10140_o_0),
    .C(n_10085_o_0),
    .Y(n_10268_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10269 (.A1(n_10061_o_0),
    .A2(n_10232_o_0),
    .B(n_10268_o_0),
    .C(n_10150_o_0),
    .Y(n_10269_o_0));
 OAI31xp33_ASAP7_75t_R n_1027 (.A1(n_878_o_0),
    .A2(n_1025_o_0),
    .A3(n_994_o_0),
    .B(n_1026_o_0),
    .Y(n_1027_o_0));
 INVx1_ASAP7_75t_R n_10270 (.A(n_10269_o_0),
    .Y(n_10270_o_0));
 OAI211xp5_ASAP7_75t_R n_10271 (.A1(n_10149_o_0),
    .A2(n_10267_o_0),
    .B(n_10270_o_0),
    .C(n_10116_o_0),
    .Y(n_10271_o_0));
 OAI31xp33_ASAP7_75t_R n_10272 (.A1(n_10067_o_0),
    .A2(n_10262_o_0),
    .A3(n_10266_o_0),
    .B(n_10271_o_0),
    .Y(n_10272_o_0));
 INVx1_ASAP7_75t_R n_10273 (.A(n_10182_o_0),
    .Y(n_10273_o_0));
 AOI22xp33_ASAP7_75t_R n_10274 (.A1(n_10273_o_0),
    .A2(n_10085_o_0),
    .B1(n_10077_o_0),
    .B2(n_10118_o_0),
    .Y(n_10274_o_0));
 OAI21xp33_ASAP7_75t_R n_10275 (.A1(n_10155_o_0),
    .A2(n_10153_o_0),
    .B(n_10177_o_0),
    .Y(n_10275_o_0));
 OAI31xp33_ASAP7_75t_R n_10276 (.A1(net56),
    .A2(n_10061_o_0),
    .A3(n_10025_o_0),
    .B(n_10275_o_0),
    .Y(n_10276_o_0));
 AOI21xp33_ASAP7_75t_R n_10277 (.A1(n_10005_o_0),
    .A2(n_10276_o_0),
    .B(n_10093_o_0),
    .Y(n_10277_o_0));
 OAI21xp33_ASAP7_75t_R n_10278 (.A1(n_10150_o_0),
    .A2(n_10274_o_0),
    .B(n_10277_o_0),
    .Y(n_10278_o_0));
 OAI21xp33_ASAP7_75t_R n_10279 (.A1(n_10040_o_0),
    .A2(n_10058_o_0),
    .B(n_10061_o_0),
    .Y(n_10279_o_0));
 NOR2xp33_ASAP7_75t_R n_1028 (.A(n_878_o_0),
    .B(n_989_o_0),
    .Y(n_1028_o_0));
 OAI31xp33_ASAP7_75t_R n_10280 (.A1(net61),
    .A2(n_10058_o_0),
    .A3(n_10043_o_0),
    .B(n_10171_o_0),
    .Y(n_10280_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10281 (.A1(n_10024_o_0),
    .A2(n_10199_o_0),
    .B(n_10279_o_0),
    .C(n_10280_o_0),
    .Y(n_10281_o_0));
 NAND3xp33_ASAP7_75t_R n_10282 (.A(n_10024_o_0),
    .B(n_10056_o_0),
    .C(net56),
    .Y(n_10282_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10283 (.A1(net24),
    .A2(n_10058_o_0),
    .B(n_10043_o_0),
    .C(n_10061_o_0),
    .Y(n_10283_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10284 (.A1(n_10282_o_0),
    .A2(n_10283_o_0),
    .B(n_10005_o_0),
    .C(n_10093_o_0),
    .Y(n_10284_o_0));
 AO21x1_ASAP7_75t_R n_10285 (.A1(n_10281_o_0),
    .A2(n_10150_o_0),
    .B(n_10284_o_0),
    .Y(n_10285_o_0));
 AOI31xp33_ASAP7_75t_R n_10286 (.A1(n_9997_o_0),
    .A2(n_10278_o_0),
    .A3(n_10285_o_0),
    .B(n_10102_o_0),
    .Y(n_10286_o_0));
 INVx1_ASAP7_75t_R n_10287 (.A(n_10188_o_0),
    .Y(n_10287_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10288 (.A1(n_10012_o_0),
    .A2(n_10043_o_0),
    .B(n_10058_o_0),
    .C(n_10077_o_0),
    .Y(n_10288_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10289 (.A1(n_10024_o_0),
    .A2(net56),
    .B(n_10288_o_0),
    .C(n_10086_o_0),
    .Y(n_10289_o_0));
 NAND2xp33_ASAP7_75t_R n_1029 (.A(n_836_o_0),
    .B(n_935_o_0),
    .Y(n_1029_o_0));
 NAND2xp33_ASAP7_75t_R n_10290 (.A(n_10012_o_0),
    .B(n_10024_o_0),
    .Y(n_10290_o_0));
 OAI211xp5_ASAP7_75t_R n_10291 (.A1(n_10037_o_0),
    .A2(n_10290_o_0),
    .B(n_10082_o_0),
    .C(n_10077_o_0),
    .Y(n_10291_o_0));
 OAI211xp5_ASAP7_75t_R n_10292 (.A1(net61),
    .A2(net56),
    .B(n_10084_o_0),
    .C(n_10085_o_0),
    .Y(n_10292_o_0));
 AOI31xp33_ASAP7_75t_R n_10293 (.A1(n_10291_o_0),
    .A2(n_10292_o_0),
    .A3(n_10146_o_0),
    .B(n_10150_o_0),
    .Y(n_10293_o_0));
 OAI21xp33_ASAP7_75t_R n_10294 (.A1(n_10093_o_0),
    .A2(n_10289_o_0),
    .B(n_10293_o_0),
    .Y(n_10294_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10295 (.A1(net56),
    .A2(n_10043_o_0),
    .B(net61),
    .C(n_10077_o_0),
    .D(n_10116_o_0),
    .Y(n_10295_o_0));
 INVx1_ASAP7_75t_R n_10296 (.A(n_10295_o_0),
    .Y(n_10296_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10297 (.A1(net24),
    .A2(net56),
    .B(n_10043_o_0),
    .C(n_10056_o_0),
    .Y(n_10297_o_0));
 OAI21xp33_ASAP7_75t_R n_10298 (.A1(n_10024_o_0),
    .A2(net61),
    .B(n_10141_o_0),
    .Y(n_10298_o_0));
 AOI21xp33_ASAP7_75t_R n_10299 (.A1(n_10159_o_0),
    .A2(n_10162_o_0),
    .B(n_10146_o_0),
    .Y(n_10299_o_0));
 NOR2xp33_ASAP7_75t_R n_1030 (.A(n_877_o_0),
    .B(n_1029_o_0),
    .Y(n_1030_o_0));
 AOI21xp33_ASAP7_75t_R n_10300 (.A1(n_10298_o_0),
    .A2(n_10299_o_0),
    .B(n_10004_o_0),
    .Y(n_10300_o_0));
 OAI21xp33_ASAP7_75t_R n_10301 (.A1(n_10296_o_0),
    .A2(n_10297_o_0),
    .B(n_10300_o_0),
    .Y(n_10301_o_0));
 OAI211xp5_ASAP7_75t_R n_10302 (.A1(n_10087_o_0),
    .A2(n_10058_o_0),
    .B(n_10077_o_0),
    .C(n_10125_o_0),
    .Y(n_10302_o_0));
 OAI211xp5_ASAP7_75t_R n_10303 (.A1(net56),
    .A2(net61),
    .B(n_10178_o_0),
    .C(n_10061_o_0),
    .Y(n_10303_o_0));
 OAI211xp5_ASAP7_75t_R n_10304 (.A1(n_10134_o_0),
    .A2(n_10043_o_0),
    .B(n_10251_o_0),
    .C(n_10061_o_0),
    .Y(n_10304_o_0));
 AOI21xp33_ASAP7_75t_R n_10305 (.A1(n_10128_o_0),
    .A2(n_10304_o_0),
    .B(n_10093_o_0),
    .Y(n_10305_o_0));
 AOI31xp33_ASAP7_75t_R n_10306 (.A1(n_10302_o_0),
    .A2(n_10303_o_0),
    .A3(n_10146_o_0),
    .B(n_10305_o_0),
    .Y(n_10306_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10307 (.A1(n_10089_o_0),
    .A2(net56),
    .B(n_10166_o_0),
    .C(n_10085_o_0),
    .Y(n_10307_o_0));
 NAND2xp33_ASAP7_75t_R n_10308 (.A(n_10149_o_0),
    .B(n_10116_o_0),
    .Y(n_10308_o_0));
 AOI21xp33_ASAP7_75t_R n_10309 (.A1(n_10012_o_0),
    .A2(n_10024_o_0),
    .B(n_10037_o_0),
    .Y(n_10309_o_0));
 AOI21xp33_ASAP7_75t_R n_1031 (.A1(n_909_o_0),
    .A2(n_1028_o_0),
    .B(n_1030_o_0),
    .Y(n_1031_o_0));
 OAI211xp5_ASAP7_75t_R n_10310 (.A1(n_10246_o_0),
    .A2(n_10309_o_0),
    .B(n_10283_o_0),
    .C(n_10149_o_0),
    .Y(n_10310_o_0));
 AOI32xp33_ASAP7_75t_R n_10311 (.A1(n_10067_o_0),
    .A2(n_10307_o_0),
    .A3(n_10078_o_0),
    .B1(n_10308_o_0),
    .B2(n_10310_o_0),
    .Y(n_10311_o_0));
 AOI21xp33_ASAP7_75t_R n_10312 (.A1(n_10306_o_0),
    .A2(n_10005_o_0),
    .B(n_10311_o_0),
    .Y(n_10312_o_0));
 INVx1_ASAP7_75t_R n_10313 (.A(n_10224_o_0),
    .Y(n_10313_o_0));
 AOI321xp33_ASAP7_75t_R n_10314 (.A1(n_10287_o_0),
    .A2(n_10294_o_0),
    .A3(n_10301_o_0),
    .B1(n_10312_o_0),
    .B2(n_9997_o_0),
    .C(n_10313_o_0),
    .Y(n_10314_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10315 (.A1(n_10188_o_0),
    .A2(n_10272_o_0),
    .B(n_10286_o_0),
    .C(n_10314_o_0),
    .Y(n_10315_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10316 (.A1(n_10106_o_0),
    .A2(n_10075_o_0),
    .B(n_10058_o_0),
    .C(n_10056_o_0),
    .Y(n_10316_o_0));
 OAI22xp33_ASAP7_75t_R n_10317 (.A1(n_10316_o_0),
    .A2(n_10245_o_0),
    .B1(n_10279_o_0),
    .B2(n_10309_o_0),
    .Y(n_10317_o_0));
 INVx1_ASAP7_75t_R n_10318 (.A(n_10317_o_0),
    .Y(n_10318_o_0));
 NAND3xp33_ASAP7_75t_R n_10319 (.A(n_10037_o_0),
    .B(n_10043_o_0),
    .C(net24),
    .Y(n_10319_o_0));
 OAI21xp33_ASAP7_75t_R n_1032 (.A1(net42),
    .A2(n_1031_o_0),
    .B(n_904_o_0),
    .Y(n_1032_o_0));
 AOI21xp33_ASAP7_75t_R n_10320 (.A1(n_10061_o_0),
    .A2(n_10319_o_0),
    .B(n_10004_o_0),
    .Y(n_10320_o_0));
 AOI21xp33_ASAP7_75t_R n_10321 (.A1(n_10298_o_0),
    .A2(n_10320_o_0),
    .B(n_10093_o_0),
    .Y(n_10321_o_0));
 OAI21xp33_ASAP7_75t_R n_10322 (.A1(n_10150_o_0),
    .A2(n_10318_o_0),
    .B(n_10321_o_0),
    .Y(n_10322_o_0));
 NOR3xp33_ASAP7_75t_R n_10323 (.A(n_10205_o_0),
    .B(n_10085_o_0),
    .C(n_10058_o_0),
    .Y(n_10323_o_0));
 AOI21xp33_ASAP7_75t_R n_10324 (.A1(n_10073_o_0),
    .A2(n_10171_o_0),
    .B(n_10005_o_0),
    .Y(n_10324_o_0));
 OAI21xp33_ASAP7_75t_R n_10325 (.A1(n_10154_o_0),
    .A2(n_10205_o_0),
    .B(n_10324_o_0),
    .Y(n_10325_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10326 (.A1(n_10004_o_0),
    .A2(n_10323_o_0),
    .B(n_10325_o_0),
    .C(n_10116_o_0),
    .Y(n_10326_o_0));
 OAI21xp33_ASAP7_75t_R n_10327 (.A1(n_10170_o_0),
    .A2(n_10156_o_0),
    .B(n_10326_o_0),
    .Y(n_10327_o_0));
 OAI21xp33_ASAP7_75t_R n_10328 (.A1(n_10205_o_0),
    .A2(n_10154_o_0),
    .B(n_10235_o_0),
    .Y(n_10328_o_0));
 NOR2xp33_ASAP7_75t_R n_10329 (.A(n_10067_o_0),
    .B(n_10150_o_0),
    .Y(n_10329_o_0));
 INVx1_ASAP7_75t_R n_1033 (.A(n_1002_o_0),
    .Y(n_1033_o_0));
 INVx1_ASAP7_75t_R n_10330 (.A(n_10288_o_0),
    .Y(n_10330_o_0));
 INVx1_ASAP7_75t_R n_10331 (.A(n_10251_o_0),
    .Y(n_10331_o_0));
 OAI211xp5_ASAP7_75t_R n_10332 (.A1(n_10330_o_0),
    .A2(n_10331_o_0),
    .B(n_10302_o_0),
    .C(n_10067_o_0),
    .Y(n_10332_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10333 (.A1(n_10087_o_0),
    .A2(net56),
    .B(n_10077_o_0),
    .C(n_10025_o_0),
    .Y(n_10333_o_0));
 OAI31xp33_ASAP7_75t_R n_10334 (.A1(n_10037_o_0),
    .A2(n_10087_o_0),
    .A3(n_10077_o_0),
    .B(n_10156_o_0),
    .Y(n_10334_o_0));
 OAI21xp33_ASAP7_75t_R n_10335 (.A1(net61),
    .A2(n_10037_o_0),
    .B(n_10056_o_0),
    .Y(n_10335_o_0));
 AOI21xp33_ASAP7_75t_R n_10336 (.A1(n_10137_o_0),
    .A2(n_10037_o_0),
    .B(n_10335_o_0),
    .Y(n_10336_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10337 (.A1(n_10333_o_0),
    .A2(n_10334_o_0),
    .B(n_10336_o_0),
    .C(n_10146_o_0),
    .Y(n_10337_o_0));
 AOI21xp33_ASAP7_75t_R n_10338 (.A1(n_10332_o_0),
    .A2(n_10337_o_0),
    .B(n_10149_o_0),
    .Y(n_10338_o_0));
 INVx1_ASAP7_75t_R n_10339 (.A(n_10141_o_0),
    .Y(n_10339_o_0));
 AOI211xp5_ASAP7_75t_R n_1034 (.A1(n_957_o_0),
    .A2(n_881_o_0),
    .B(n_892_o_0),
    .C(n_877_o_0),
    .Y(n_1034_o_0));
 OAI22xp33_ASAP7_75t_R n_10340 (.A1(n_10107_o_0),
    .A2(n_10261_o_0),
    .B1(n_10339_o_0),
    .B2(n_10111_o_0),
    .Y(n_10340_o_0));
 OAI21xp33_ASAP7_75t_R n_10341 (.A1(n_10308_o_0),
    .A2(n_10340_o_0),
    .B(n_10313_o_0),
    .Y(n_10341_o_0));
 AOI211xp5_ASAP7_75t_R n_10342 (.A1(n_10328_o_0),
    .A2(n_10329_o_0),
    .B(n_10338_o_0),
    .C(n_10341_o_0),
    .Y(n_10342_o_0));
 AOI31xp33_ASAP7_75t_R n_10343 (.A1(n_10224_o_0),
    .A2(n_10322_o_0),
    .A3(n_10327_o_0),
    .B(n_10342_o_0),
    .Y(n_10343_o_0));
 AOI31xp33_ASAP7_75t_R n_10344 (.A1(n_10085_o_0),
    .A2(n_10112_o_0),
    .A3(n_10143_o_0),
    .B(n_10116_o_0),
    .Y(n_10344_o_0));
 OAI21xp33_ASAP7_75t_R n_10345 (.A1(n_10037_o_0),
    .A2(n_10068_o_0),
    .B(n_10135_o_0),
    .Y(n_10345_o_0));
 OAI221xp5_ASAP7_75t_R n_10346 (.A1(net61),
    .A2(n_10043_o_0),
    .B1(n_10037_o_0),
    .B2(n_10075_o_0),
    .C(n_10077_o_0),
    .Y(n_10346_o_0));
 OAI211xp5_ASAP7_75t_R n_10347 (.A1(n_10137_o_0),
    .A2(net56),
    .B(n_10118_o_0),
    .C(n_10085_o_0),
    .Y(n_10347_o_0));
 AOI21xp33_ASAP7_75t_R n_10348 (.A1(n_10346_o_0),
    .A2(n_10347_o_0),
    .B(n_10146_o_0),
    .Y(n_10348_o_0));
 AOI21xp33_ASAP7_75t_R n_10349 (.A1(n_10344_o_0),
    .A2(n_10345_o_0),
    .B(n_10348_o_0),
    .Y(n_10349_o_0));
 OAI21xp33_ASAP7_75t_R n_1035 (.A1(n_877_o_0),
    .A2(n_886_o_0),
    .B(n_829_o_0),
    .Y(n_1035_o_0));
 NOR2xp33_ASAP7_75t_R n_10350 (.A(n_10037_o_0),
    .B(n_10068_o_0),
    .Y(n_10350_o_0));
 AOI211xp5_ASAP7_75t_R n_10351 (.A1(n_10205_o_0),
    .A2(n_10037_o_0),
    .B(n_10061_o_0),
    .C(n_10350_o_0),
    .Y(n_10351_o_0));
 NAND3xp33_ASAP7_75t_R n_10352 (.A(n_10170_o_0),
    .B(n_10134_o_0),
    .C(n_10140_o_0),
    .Y(n_10352_o_0));
 OAI32xp33_ASAP7_75t_R n_10353 (.A1(n_10116_o_0),
    .A2(n_10351_o_0),
    .A3(n_10226_o_0),
    .B1(n_10093_o_0),
    .B2(n_10352_o_0),
    .Y(n_10353_o_0));
 OAI22xp33_ASAP7_75t_R n_10354 (.A1(n_10349_o_0),
    .A2(n_10004_o_0),
    .B1(n_10353_o_0),
    .B2(n_10150_o_0),
    .Y(n_10354_o_0));
 OAI21xp33_ASAP7_75t_R n_10355 (.A1(n_10151_o_0),
    .A2(n_10176_o_0),
    .B(n_10249_o_0),
    .Y(n_10355_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10356 (.A1(n_10068_o_0),
    .A2(n_10037_o_0),
    .B(n_10245_o_0),
    .C(n_10085_o_0),
    .Y(n_10356_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10357 (.A1(n_10309_o_0),
    .A2(n_10316_o_0),
    .B(n_10356_o_0),
    .C(n_10067_o_0),
    .Y(n_10357_o_0));
 AOI21xp33_ASAP7_75t_R n_10358 (.A1(n_10116_o_0),
    .A2(n_10355_o_0),
    .B(n_10357_o_0),
    .Y(n_10358_o_0));
 AOI21xp33_ASAP7_75t_R n_10359 (.A1(net56),
    .A2(n_10137_o_0),
    .B(n_10279_o_0),
    .Y(n_10359_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1036 (.A1(n_877_o_0),
    .A2(n_953_o_0),
    .B(n_1035_o_0),
    .C(n_903_o_0),
    .Y(n_1036_o_0));
 OAI211xp5_ASAP7_75t_R n_10360 (.A1(n_10280_o_0),
    .A2(n_10093_o_0),
    .B(n_10149_o_0),
    .C(n_10296_o_0),
    .Y(n_10360_o_0));
 AOI211xp5_ASAP7_75t_R n_10361 (.A1(n_10116_o_0),
    .A2(n_10359_o_0),
    .B(n_10360_o_0),
    .C(n_10188_o_0),
    .Y(n_10361_o_0));
 AOI211xp5_ASAP7_75t_R n_10362 (.A1(n_10358_o_0),
    .A2(n_10150_o_0),
    .B(n_10361_o_0),
    .C(n_10313_o_0),
    .Y(n_10362_o_0));
 AOI211xp5_ASAP7_75t_R n_10363 (.A1(net61),
    .A2(n_10043_o_0),
    .B(n_10263_o_0),
    .C(n_10061_o_0),
    .Y(n_10363_o_0));
 AOI21xp33_ASAP7_75t_R n_10364 (.A1(n_10124_o_0),
    .A2(n_10091_o_0),
    .B(n_10363_o_0),
    .Y(n_10364_o_0));
 INVx1_ASAP7_75t_R n_10365 (.A(n_10309_o_0),
    .Y(n_10365_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10366 (.A1(net24),
    .A2(n_10037_o_0),
    .B(n_10319_o_0),
    .C(n_10056_o_0),
    .Y(n_10366_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10367 (.A1(n_10365_o_0),
    .A2(n_10135_o_0),
    .B(n_10366_o_0),
    .C(n_10093_o_0),
    .Y(n_10367_o_0));
 OAI21xp33_ASAP7_75t_R n_10368 (.A1(n_10146_o_0),
    .A2(n_10364_o_0),
    .B(n_10367_o_0),
    .Y(n_10368_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10369 (.A1(n_10149_o_0),
    .A2(n_10368_o_0),
    .B(n_10224_o_0),
    .C(n_10287_o_0),
    .Y(n_10369_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1037 (.A1(n_1033_o_0),
    .A2(n_1034_o_0),
    .B(n_891_o_0),
    .C(n_1036_o_0),
    .Y(n_1037_o_0));
 AOI211xp5_ASAP7_75t_R n_10370 (.A1(n_10354_o_0),
    .A2(n_10103_o_0),
    .B(n_10362_o_0),
    .C(n_10369_o_0),
    .Y(n_10370_o_0));
 AOI21xp33_ASAP7_75t_R n_10371 (.A1(n_9997_o_0),
    .A2(n_10343_o_0),
    .B(n_10370_o_0),
    .Y(n_10371_o_0));
 AOI21xp33_ASAP7_75t_R n_10372 (.A1(net56),
    .A2(n_10024_o_0),
    .B(n_10061_o_0),
    .Y(n_10372_o_0));
 NAND2xp33_ASAP7_75t_R n_10373 (.A(n_10085_o_0),
    .B(n_10125_o_0),
    .Y(n_10373_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10374 (.A1(n_10037_o_0),
    .A2(n_10089_o_0),
    .B(n_10373_o_0),
    .C(n_10146_o_0),
    .Y(n_10374_o_0));
 AOI21xp33_ASAP7_75t_R n_10375 (.A1(n_10124_o_0),
    .A2(n_10372_o_0),
    .B(n_10374_o_0),
    .Y(n_10375_o_0));
 OAI21xp33_ASAP7_75t_R n_10376 (.A1(n_10109_o_0),
    .A2(n_10339_o_0),
    .B(n_10067_o_0),
    .Y(n_10376_o_0));
 AOI21xp33_ASAP7_75t_R n_10377 (.A1(net56),
    .A2(n_10085_o_0),
    .B(n_10376_o_0),
    .Y(n_10377_o_0));
 AOI31xp33_ASAP7_75t_R n_10378 (.A1(n_10077_o_0),
    .A2(n_10076_o_0),
    .A3(n_10119_o_0),
    .B(n_10093_o_0),
    .Y(n_10378_o_0));
 INVx1_ASAP7_75t_R n_10379 (.A(n_10378_o_0),
    .Y(n_10379_o_0));
 AOI21xp33_ASAP7_75t_R n_1038 (.A1(n_985_o_0),
    .A2(n_1037_o_0),
    .B(n_931_o_0),
    .Y(n_1038_o_0));
 INVx1_ASAP7_75t_R n_10380 (.A(n_10206_o_0),
    .Y(n_10380_o_0));
 AOI21xp33_ASAP7_75t_R n_10381 (.A1(n_10058_o_0),
    .A2(n_10156_o_0),
    .B(n_10061_o_0),
    .Y(n_10381_o_0));
 AOI21xp33_ASAP7_75t_R n_10382 (.A1(n_10085_o_0),
    .A2(n_10380_o_0),
    .B(n_10381_o_0),
    .Y(n_10382_o_0));
 AOI21xp33_ASAP7_75t_R n_10383 (.A1(n_10146_o_0),
    .A2(n_10382_o_0),
    .B(n_10004_o_0),
    .Y(n_10383_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10384 (.A1(n_10092_o_0),
    .A2(n_10091_o_0),
    .B(n_10379_o_0),
    .C(n_10383_o_0),
    .Y(n_10384_o_0));
 OAI31xp33_ASAP7_75t_R n_10385 (.A1(n_10150_o_0),
    .A2(n_10375_o_0),
    .A3(n_10377_o_0),
    .B(n_10384_o_0),
    .Y(n_10385_o_0));
 AOI211xp5_ASAP7_75t_R n_10386 (.A1(n_10043_o_0),
    .A2(n_10037_o_0),
    .B(n_10219_o_0),
    .C(n_10061_o_0),
    .Y(n_10386_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10387 (.A1(n_10137_o_0),
    .A2(n_10037_o_0),
    .B(n_10071_o_0),
    .C(n_10386_o_0),
    .Y(n_10387_o_0));
 AOI21xp33_ASAP7_75t_R n_10388 (.A1(n_10144_o_0),
    .A2(n_10057_o_0),
    .B(n_10146_o_0),
    .Y(n_10388_o_0));
 AOI211xp5_ASAP7_75t_R n_10389 (.A1(n_10093_o_0),
    .A2(n_10387_o_0),
    .B(n_10388_o_0),
    .C(n_10005_o_0),
    .Y(n_10389_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1039 (.A1(net16),
    .A2(n_1027_o_0),
    .B(n_1032_o_0),
    .C(n_1038_o_0),
    .Y(n_1039_o_0));
 NAND2xp33_ASAP7_75t_R n_10390 (.A(n_10203_o_0),
    .B(n_10112_o_0),
    .Y(n_10390_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10391 (.A1(n_10056_o_0),
    .A2(n_10242_o_0),
    .B(n_10390_o_0),
    .C(n_10350_o_0),
    .Y(n_10391_o_0));
 NOR3xp33_ASAP7_75t_R n_10392 (.A(n_10087_o_0),
    .B(n_10077_o_0),
    .C(n_10037_o_0),
    .Y(n_10392_o_0));
 OAI21xp33_ASAP7_75t_R n_10393 (.A1(n_10085_o_0),
    .A2(n_10290_o_0),
    .B(n_10116_o_0),
    .Y(n_10393_o_0));
 OAI21xp33_ASAP7_75t_R n_10394 (.A1(n_10392_o_0),
    .A2(n_10393_o_0),
    .B(n_10150_o_0),
    .Y(n_10394_o_0));
 AOI21xp33_ASAP7_75t_R n_10395 (.A1(n_10093_o_0),
    .A2(n_10391_o_0),
    .B(n_10394_o_0),
    .Y(n_10395_o_0));
 OAI21xp33_ASAP7_75t_R n_10396 (.A1(n_10389_o_0),
    .A2(n_10395_o_0),
    .B(n_9997_o_0),
    .Y(n_10396_o_0));
 OAI21xp33_ASAP7_75t_R n_10397 (.A1(n_10188_o_0),
    .A2(n_10385_o_0),
    .B(n_10396_o_0),
    .Y(n_10397_o_0));
 AOI211xp5_ASAP7_75t_R n_10398 (.A1(net56),
    .A2(n_10087_o_0),
    .B(n_10331_o_0),
    .C(n_10085_o_0),
    .Y(n_10398_o_0));
 NOR2xp33_ASAP7_75t_R n_10399 (.A(n_10037_o_0),
    .B(n_10059_o_0),
    .Y(n_10399_o_0));
 OAI31xp33_ASAP7_75t_R n_1040 (.A1(n_1018_o_0),
    .A2(n_1024_o_0),
    .A3(n_930_o_0),
    .B(n_1039_o_0),
    .Y(n_1040_o_0));
 OAI321xp33_ASAP7_75t_R n_10400 (.A1(n_10166_o_0),
    .A2(n_10399_o_0),
    .A3(n_10085_o_0),
    .B1(n_10373_o_0),
    .B2(n_10151_o_0),
    .C(n_10004_o_0),
    .Y(n_10400_o_0));
 OAI31xp33_ASAP7_75t_R n_10401 (.A1(n_10004_o_0),
    .A2(n_10168_o_0),
    .A3(n_10398_o_0),
    .B(n_10400_o_0),
    .Y(n_10401_o_0));
 OAI321xp33_ASAP7_75t_R n_10402 (.A1(n_10037_o_0),
    .A2(n_10077_o_0),
    .A3(n_10087_o_0),
    .B1(n_10089_o_0),
    .B2(n_10090_o_0),
    .C(n_10082_o_0),
    .Y(n_10402_o_0));
 AOI31xp33_ASAP7_75t_R n_10403 (.A1(n_10077_o_0),
    .A2(n_10108_o_0),
    .A3(n_10119_o_0),
    .B(n_10005_o_0),
    .Y(n_10403_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10404 (.A1(n_10024_o_0),
    .A2(n_10218_o_0),
    .B(n_10373_o_0),
    .C(n_10403_o_0),
    .Y(n_10404_o_0));
 OAI211xp5_ASAP7_75t_R n_10405 (.A1(n_10402_o_0),
    .A2(n_10004_o_0),
    .B(n_10146_o_0),
    .C(n_10404_o_0),
    .Y(n_10405_o_0));
 OAI211xp5_ASAP7_75t_R n_10406 (.A1(n_10401_o_0),
    .A2(n_10093_o_0),
    .B(n_10188_o_0),
    .C(n_10405_o_0),
    .Y(n_10406_o_0));
 NAND2xp33_ASAP7_75t_R n_10407 (.A(n_10268_o_0),
    .B(n_10235_o_0),
    .Y(n_10407_o_0));
 INVx1_ASAP7_75t_R n_10408 (.A(n_10241_o_0),
    .Y(n_10408_o_0));
 OAI21xp33_ASAP7_75t_R n_10409 (.A1(n_10218_o_0),
    .A2(n_10408_o_0),
    .B(n_10237_o_0),
    .Y(n_10409_o_0));
 AOI211xp5_ASAP7_75t_R n_1041 (.A1(n_881_o_0),
    .A2(n_933_o_0),
    .B(n_877_o_0),
    .C(n_859_o_0),
    .Y(n_1041_o_0));
 OAI21xp33_ASAP7_75t_R n_10410 (.A1(n_10005_o_0),
    .A2(n_10407_o_0),
    .B(n_10409_o_0),
    .Y(n_10410_o_0));
 NAND3xp33_ASAP7_75t_R n_10411 (.A(n_10167_o_0),
    .B(n_10124_o_0),
    .C(n_10005_o_0),
    .Y(n_10411_o_0));
 OAI21xp33_ASAP7_75t_R n_10412 (.A1(n_10037_o_0),
    .A2(n_10156_o_0),
    .B(n_10085_o_0),
    .Y(n_10412_o_0));
 AOI21xp33_ASAP7_75t_R n_10413 (.A1(n_10043_o_0),
    .A2(n_10037_o_0),
    .B(n_10061_o_0),
    .Y(n_10413_o_0));
 AOI21xp33_ASAP7_75t_R n_10414 (.A1(n_10413_o_0),
    .A2(n_10225_o_0),
    .B(n_10150_o_0),
    .Y(n_10414_o_0));
 OAI21xp33_ASAP7_75t_R n_10415 (.A1(n_10412_o_0),
    .A2(n_10129_o_0),
    .B(n_10414_o_0),
    .Y(n_10415_o_0));
 AOI31xp33_ASAP7_75t_R n_10416 (.A1(n_10411_o_0),
    .A2(n_10415_o_0),
    .A3(n_10146_o_0),
    .B(n_9997_o_0),
    .Y(n_10416_o_0));
 OAI21xp33_ASAP7_75t_R n_10417 (.A1(n_10093_o_0),
    .A2(n_10410_o_0),
    .B(n_10416_o_0),
    .Y(n_10417_o_0));
 AOI21xp33_ASAP7_75t_R n_10418 (.A1(n_10406_o_0),
    .A2(n_10417_o_0),
    .B(n_10102_o_0),
    .Y(n_10418_o_0));
 AOI21xp33_ASAP7_75t_R n_10419 (.A1(n_10102_o_0),
    .A2(n_10397_o_0),
    .B(n_10418_o_0),
    .Y(n_10419_o_0));
 AOI211xp5_ASAP7_75t_R n_1042 (.A1(n_860_o_0),
    .A2(net32),
    .B(n_878_o_0),
    .C(n_907_o_0),
    .Y(n_1042_o_0));
 AOI211xp5_ASAP7_75t_R n_10420 (.A1(n_10137_o_0),
    .A2(n_10058_o_0),
    .B(n_10166_o_0),
    .C(n_10085_o_0),
    .Y(n_10420_o_0));
 AOI211xp5_ASAP7_75t_R n_10421 (.A1(net61),
    .A2(n_10288_o_0),
    .B(n_10420_o_0),
    .C(n_10067_o_0),
    .Y(n_10421_o_0));
 OAI211xp5_ASAP7_75t_R n_10422 (.A1(n_10062_o_0),
    .A2(n_10309_o_0),
    .B(n_10126_o_0),
    .C(n_10116_o_0),
    .Y(n_10422_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10423 (.A1(n_10092_o_0),
    .A2(n_10069_o_0),
    .B(n_10056_o_0),
    .C(n_10146_o_0),
    .Y(n_10423_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10424 (.A1(n_10085_o_0),
    .A2(n_10024_o_0),
    .B(n_10386_o_0),
    .C(n_10067_o_0),
    .Y(n_10424_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10425 (.A1(n_10225_o_0),
    .A2(n_10120_o_0),
    .B(n_10423_o_0),
    .C(n_10424_o_0),
    .Y(n_10425_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10426 (.A1(n_9990_o_0),
    .A2(n_9995_o_0),
    .B(n_9996_o_0),
    .C(n_10421_o_0),
    .Y(n_10426_o_0));
 OAI321xp33_ASAP7_75t_R n_10427 (.A1(n_10421_o_0),
    .A2(n_10422_o_0),
    .A3(n_9997_o_0),
    .B1(n_10287_o_0),
    .B2(n_10425_o_0),
    .C(n_10426_o_0),
    .Y(n_10427_o_0));
 OAI21xp33_ASAP7_75t_R n_10428 (.A1(n_10037_o_0),
    .A2(n_10111_o_0),
    .B(n_10146_o_0),
    .Y(n_10428_o_0));
 AOI21xp33_ASAP7_75t_R n_10429 (.A1(n_10077_o_0),
    .A2(n_10119_o_0),
    .B(n_10428_o_0),
    .Y(n_10429_o_0));
 AOI31xp33_ASAP7_75t_R n_1043 (.A1(n_933_o_0),
    .A2(net32),
    .A3(n_877_o_0),
    .B(n_891_o_0),
    .Y(n_1043_o_0));
 AOI31xp33_ASAP7_75t_R n_10430 (.A1(n_10116_o_0),
    .A2(n_10316_o_0),
    .A3(n_10356_o_0),
    .B(n_10429_o_0),
    .Y(n_10430_o_0));
 AOI211xp5_ASAP7_75t_R n_10431 (.A1(net24),
    .A2(net56),
    .B(n_10024_o_0),
    .C(n_10061_o_0),
    .Y(n_10431_o_0));
 AOI31xp33_ASAP7_75t_R n_10432 (.A1(n_10085_o_0),
    .A2(n_10205_o_0),
    .A3(net56),
    .B(n_10431_o_0),
    .Y(n_10432_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10433 (.A1(n_10037_o_0),
    .A2(n_10290_o_0),
    .B(n_10056_o_0),
    .C(n_10146_o_0),
    .Y(n_10433_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10434 (.A1(n_10044_o_0),
    .A2(n_10107_o_0),
    .B(n_10433_o_0),
    .C(n_10257_o_0),
    .Y(n_10434_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10435 (.A1(n_10067_o_0),
    .A2(n_10432_o_0),
    .B(n_10434_o_0),
    .C(n_10150_o_0),
    .Y(n_10435_o_0));
 OAI21xp33_ASAP7_75t_R n_10436 (.A1(n_10188_o_0),
    .A2(n_10430_o_0),
    .B(n_10435_o_0),
    .Y(n_10436_o_0));
 OA21x2_ASAP7_75t_R n_10437 (.A1(n_10427_o_0),
    .A2(n_10004_o_0),
    .B(n_10436_o_0),
    .Y(n_10437_o_0));
 OAI21xp33_ASAP7_75t_R n_10438 (.A1(n_10155_o_0),
    .A2(n_10153_o_0),
    .B(n_10118_o_0),
    .Y(n_10438_o_0));
 OAI31xp33_ASAP7_75t_R n_10439 (.A1(n_10061_o_0),
    .A2(n_10242_o_0),
    .A3(n_10350_o_0),
    .B(n_10438_o_0),
    .Y(n_10439_o_0));
 INVx1_ASAP7_75t_R n_1044 (.A(n_889_o_0),
    .Y(n_1044_o_0));
 NAND3xp33_ASAP7_75t_R n_10440 (.A(n_10137_o_0),
    .B(n_10085_o_0),
    .C(net56),
    .Y(n_10440_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10441 (.A1(n_10061_o_0),
    .A2(n_10109_o_0),
    .B(n_10440_o_0),
    .C(n_10194_o_0),
    .Y(n_10441_o_0));
 AOI22xp33_ASAP7_75t_R n_10442 (.A1(n_10439_o_0),
    .A2(n_10005_o_0),
    .B1(n_10149_o_0),
    .B2(n_10441_o_0),
    .Y(n_10442_o_0));
 NAND2xp33_ASAP7_75t_R n_10443 (.A(n_10177_o_0),
    .B(n_10110_o_0),
    .Y(n_10443_o_0));
 OAI31xp33_ASAP7_75t_R n_10444 (.A1(n_10056_o_0),
    .A2(n_10194_o_0),
    .A3(n_10195_o_0),
    .B(n_10443_o_0),
    .Y(n_10444_o_0));
 NAND2xp33_ASAP7_75t_R n_10445 (.A(n_10116_o_0),
    .B(n_10005_o_0),
    .Y(n_10445_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10446 (.A1(net61),
    .A2(n_10056_o_0),
    .B(n_10142_o_0),
    .C(n_10445_o_0),
    .Y(n_10446_o_0));
 AOI31xp33_ASAP7_75t_R n_10447 (.A1(n_10116_o_0),
    .A2(n_10149_o_0),
    .A3(n_10444_o_0),
    .B(n_10446_o_0),
    .Y(n_10447_o_0));
 OAI21xp33_ASAP7_75t_R n_10448 (.A1(n_10067_o_0),
    .A2(n_10442_o_0),
    .B(n_10447_o_0),
    .Y(n_10448_o_0));
 NOR2xp33_ASAP7_75t_R n_10449 (.A(n_10058_o_0),
    .B(n_10087_o_0),
    .Y(n_10449_o_0));
 NAND3xp33_ASAP7_75t_R n_1045 (.A(n_1044_o_0),
    .B(net32),
    .C(n_878_o_0),
    .Y(n_1045_o_0));
 OAI21xp33_ASAP7_75t_R n_10450 (.A1(n_10155_o_0),
    .A2(n_10153_o_0),
    .B(n_10069_o_0),
    .Y(n_10450_o_0));
 OAI31xp33_ASAP7_75t_R n_10451 (.A1(n_10061_o_0),
    .A2(n_10109_o_0),
    .A3(n_10449_o_0),
    .B(n_10450_o_0),
    .Y(n_10451_o_0));
 AOI31xp33_ASAP7_75t_R n_10452 (.A1(net56),
    .A2(n_10059_o_0),
    .A3(n_10056_o_0),
    .B(n_10004_o_0),
    .Y(n_10452_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10453 (.A1(n_10077_o_0),
    .A2(n_10309_o_0),
    .B(n_10452_o_0),
    .C(n_10067_o_0),
    .Y(n_10453_o_0));
 OAI21xp33_ASAP7_75t_R n_10454 (.A1(n_10005_o_0),
    .A2(n_10451_o_0),
    .B(n_10453_o_0),
    .Y(n_10454_o_0));
 NAND2xp33_ASAP7_75t_R n_10455 (.A(n_10279_o_0),
    .B(n_10005_o_0),
    .Y(n_10455_o_0));
 AND3x1_ASAP7_75t_R n_10456 (.A(n_10092_o_0),
    .B(n_10118_o_0),
    .C(n_10077_o_0),
    .Y(n_10456_o_0));
 AOI21xp33_ASAP7_75t_R n_10457 (.A1(n_10137_o_0),
    .A2(n_10085_o_0),
    .B(n_10005_o_0),
    .Y(n_10457_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10458 (.A1(n_10061_o_0),
    .A2(n_10194_o_0),
    .B(n_10457_o_0),
    .C(n_10146_o_0),
    .Y(n_10458_o_0));
 OAI21xp33_ASAP7_75t_R n_10459 (.A1(n_10455_o_0),
    .A2(n_10456_o_0),
    .B(n_10458_o_0),
    .Y(n_10459_o_0));
 NAND2xp33_ASAP7_75t_R n_1046 (.A(n_878_o_0),
    .B(n_861_o_0),
    .Y(n_1046_o_0));
 AOI31xp33_ASAP7_75t_R n_10460 (.A1(n_9997_o_0),
    .A2(n_10454_o_0),
    .A3(n_10459_o_0),
    .B(n_10313_o_0),
    .Y(n_10460_o_0));
 OAI21xp33_ASAP7_75t_R n_10461 (.A1(n_10188_o_0),
    .A2(n_10448_o_0),
    .B(n_10460_o_0),
    .Y(n_10461_o_0));
 OAI21xp33_ASAP7_75t_R n_10462 (.A1(n_10102_o_0),
    .A2(n_10437_o_0),
    .B(n_10461_o_0),
    .Y(n_10462_o_0));
 NAND3xp33_ASAP7_75t_R n_10463 (.A(n_10112_o_0),
    .B(n_10125_o_0),
    .C(n_10085_o_0),
    .Y(n_10463_o_0));
 OAI211xp5_ASAP7_75t_R n_10464 (.A1(n_10024_o_0),
    .A2(n_10085_o_0),
    .B(n_10463_o_0),
    .C(n_10150_o_0),
    .Y(n_10464_o_0));
 NAND3xp33_ASAP7_75t_R n_10465 (.A(n_10124_o_0),
    .B(n_10127_o_0),
    .C(n_10125_o_0),
    .Y(n_10465_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10466 (.A1(n_10137_o_0),
    .A2(net56),
    .B(n_10208_o_0),
    .C(n_10149_o_0),
    .Y(n_10466_o_0));
 AO21x1_ASAP7_75t_R n_10467 (.A1(n_10465_o_0),
    .A2(n_10061_o_0),
    .B(n_10466_o_0),
    .Y(n_10467_o_0));
 AO21x1_ASAP7_75t_R n_10468 (.A1(n_10464_o_0),
    .A2(n_10467_o_0),
    .B(n_10093_o_0),
    .Y(n_10468_o_0));
 OAI21xp33_ASAP7_75t_R n_10469 (.A1(net24),
    .A2(n_10154_o_0),
    .B(n_10004_o_0),
    .Y(n_10469_o_0));
 NAND4xp25_ASAP7_75t_R n_1047 (.A(n_1043_o_0),
    .B(n_1045_o_0),
    .C(n_975_o_0),
    .D(n_1046_o_0),
    .Y(n_1047_o_0));
 AO21x1_ASAP7_75t_R n_10470 (.A1(n_10076_o_0),
    .A2(n_10141_o_0),
    .B(n_10469_o_0),
    .Y(n_10470_o_0));
 OAI21xp33_ASAP7_75t_R n_10471 (.A1(n_10056_o_0),
    .A2(n_10178_o_0),
    .B(n_10150_o_0),
    .Y(n_10471_o_0));
 AO21x1_ASAP7_75t_R n_10472 (.A1(n_10203_o_0),
    .A2(n_10156_o_0),
    .B(n_10471_o_0),
    .Y(n_10472_o_0));
 AOI21xp33_ASAP7_75t_R n_10473 (.A1(n_10470_o_0),
    .A2(n_10472_o_0),
    .B(n_10116_o_0),
    .Y(n_10473_o_0));
 OAI21xp33_ASAP7_75t_R n_10474 (.A1(n_10319_o_0),
    .A2(n_10056_o_0),
    .B(n_10473_o_0),
    .Y(n_10474_o_0));
 AOI211xp5_ASAP7_75t_R n_10475 (.A1(n_10156_o_0),
    .A2(net56),
    .B(n_10449_o_0),
    .C(n_10061_o_0),
    .Y(n_10475_o_0));
 AOI211xp5_ASAP7_75t_R n_10476 (.A1(n_10195_o_0),
    .A2(n_10024_o_0),
    .B(n_10056_o_0),
    .C(n_10242_o_0),
    .Y(n_10476_o_0));
 NAND2xp33_ASAP7_75t_R n_10477 (.A(n_10085_o_0),
    .B(n_10172_o_0),
    .Y(n_10477_o_0));
 OAI211xp5_ASAP7_75t_R n_10478 (.A1(n_10025_o_0),
    .A2(n_10119_o_0),
    .B(n_10077_o_0),
    .C(n_10076_o_0),
    .Y(n_10478_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10479 (.A1(net24),
    .A2(net56),
    .B(n_10477_o_0),
    .C(n_10478_o_0),
    .Y(n_10479_o_0));
 OAI311xp33_ASAP7_75t_R n_1048 (.A1(net16),
    .A2(n_1041_o_0),
    .A3(n_1042_o_0),
    .B1(n_904_o_0),
    .C1(n_1047_o_0),
    .Y(n_1048_o_0));
 OAI32xp33_ASAP7_75t_R n_10480 (.A1(n_10149_o_0),
    .A2(n_10475_o_0),
    .A3(n_10476_o_0),
    .B1(n_10479_o_0),
    .B2(n_10005_o_0),
    .Y(n_10480_o_0));
 NOR2xp33_ASAP7_75t_R n_10481 (.A(net61),
    .B(n_10058_o_0),
    .Y(n_10481_o_0));
 OAI21xp33_ASAP7_75t_R n_10482 (.A1(n_10037_o_0),
    .A2(n_10068_o_0),
    .B(n_10056_o_0),
    .Y(n_10482_o_0));
 OAI311xp33_ASAP7_75t_R n_10483 (.A1(n_10043_o_0),
    .A2(n_10056_o_0),
    .A3(n_10481_o_0),
    .B1(n_10149_o_0),
    .C1(n_10482_o_0),
    .Y(n_10483_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10484 (.A1(n_10004_o_0),
    .A2(n_10274_o_0),
    .B(n_10483_o_0),
    .C(n_10323_o_0),
    .Y(n_10484_o_0));
 AOI21xp33_ASAP7_75t_R n_10485 (.A1(n_10093_o_0),
    .A2(n_10484_o_0),
    .B(n_10257_o_0),
    .Y(n_10485_o_0));
 OAI21xp33_ASAP7_75t_R n_10486 (.A1(n_10146_o_0),
    .A2(n_10480_o_0),
    .B(n_10485_o_0),
    .Y(n_10486_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10487 (.A1(n_10468_o_0),
    .A2(n_10474_o_0),
    .B(n_10188_o_0),
    .C(n_10486_o_0),
    .Y(n_10487_o_0));
 AOI21xp33_ASAP7_75t_R n_10488 (.A1(n_10024_o_0),
    .A2(net56),
    .B(n_10129_o_0),
    .Y(n_10488_o_0));
 INVx1_ASAP7_75t_R n_10489 (.A(n_10413_o_0),
    .Y(n_10489_o_0));
 OAI31xp33_ASAP7_75t_R n_1049 (.A1(n_878_o_0),
    .A2(n_915_o_0),
    .A3(n_949_o_0),
    .B(n_1013_o_0),
    .Y(n_1049_o_0));
 OAI22xp33_ASAP7_75t_R n_10490 (.A1(n_10488_o_0),
    .A2(n_10056_o_0),
    .B1(n_10350_o_0),
    .B2(n_10489_o_0),
    .Y(n_10490_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10491 (.A1(net24),
    .A2(net56),
    .B(n_10085_o_0),
    .C(n_10093_o_0),
    .Y(n_10491_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10492 (.A1(n_10037_o_0),
    .A2(n_10290_o_0),
    .B(n_10088_o_0),
    .C(n_10491_o_0),
    .Y(n_10492_o_0));
 AOI21xp33_ASAP7_75t_R n_10493 (.A1(n_10116_o_0),
    .A2(n_10490_o_0),
    .B(n_10492_o_0),
    .Y(n_10493_o_0));
 OAI21xp33_ASAP7_75t_R n_10494 (.A1(n_10037_o_0),
    .A2(n_10137_o_0),
    .B(n_10056_o_0),
    .Y(n_10494_o_0));
 OAI211xp5_ASAP7_75t_R n_10495 (.A1(n_10129_o_0),
    .A2(n_10167_o_0),
    .B(n_10329_o_0),
    .C(n_10494_o_0),
    .Y(n_10495_o_0));
 OAI21xp33_ASAP7_75t_R n_10496 (.A1(n_10308_o_0),
    .A2(n_10307_o_0),
    .B(n_10495_o_0),
    .Y(n_10496_o_0));
 AOI21xp33_ASAP7_75t_R n_10497 (.A1(n_10005_o_0),
    .A2(n_10493_o_0),
    .B(n_10496_o_0),
    .Y(n_10497_o_0));
 INVx1_ASAP7_75t_R n_10498 (.A(n_10117_o_0),
    .Y(n_10498_o_0));
 OAI211xp5_ASAP7_75t_R n_10499 (.A1(n_10159_o_0),
    .A2(n_10061_o_0),
    .B(n_10356_o_0),
    .C(n_10067_o_0),
    .Y(n_10499_o_0));
 INVx1_ASAP7_75t_R n_1050 (.A(n_882_o_0),
    .Y(n_1050_o_0));
 OAI21xp33_ASAP7_75t_R n_10500 (.A1(n_10241_o_0),
    .A2(n_10498_o_0),
    .B(n_10499_o_0),
    .Y(n_10500_o_0));
 OAI21xp33_ASAP7_75t_R n_10501 (.A1(net24),
    .A2(n_10024_o_0),
    .B(n_10061_o_0),
    .Y(n_10501_o_0));
 AOI21xp33_ASAP7_75t_R n_10502 (.A1(n_10501_o_0),
    .A2(n_10208_o_0),
    .B(n_10199_o_0),
    .Y(n_10502_o_0));
 OAI21xp33_ASAP7_75t_R n_10503 (.A1(net61),
    .A2(n_10056_o_0),
    .B(n_10043_o_0),
    .Y(n_10503_o_0));
 AOI31xp33_ASAP7_75t_R n_10504 (.A1(n_10116_o_0),
    .A2(n_10503_o_0),
    .A3(n_10143_o_0),
    .B(n_10149_o_0),
    .Y(n_10504_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10505 (.A1(n_10067_o_0),
    .A2(n_10502_o_0),
    .B(n_10504_o_0),
    .C(n_9997_o_0),
    .Y(n_10505_o_0));
 OAI21xp33_ASAP7_75t_R n_10506 (.A1(n_10005_o_0),
    .A2(n_10500_o_0),
    .B(n_10505_o_0),
    .Y(n_10506_o_0));
 OAI21xp33_ASAP7_75t_R n_10507 (.A1(n_10287_o_0),
    .A2(n_10497_o_0),
    .B(n_10506_o_0),
    .Y(n_10507_o_0));
 OAI22xp33_ASAP7_75t_R n_10508 (.A1(n_10487_o_0),
    .A2(n_10102_o_0),
    .B1(n_10507_o_0),
    .B2(n_10313_o_0),
    .Y(n_10508_o_0));
 OAI21xp33_ASAP7_75t_R n_10509 (.A1(n_10241_o_0),
    .A2(n_10381_o_0),
    .B(n_10124_o_0),
    .Y(n_10509_o_0));
 AOI21xp33_ASAP7_75t_R n_1051 (.A1(n_881_o_0),
    .A2(n_913_o_0),
    .B(n_878_o_0),
    .Y(n_1051_o_0));
 INVx1_ASAP7_75t_R n_10510 (.A(n_10449_o_0),
    .Y(n_10510_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10511 (.A1(n_10061_o_0),
    .A2(n_10206_o_0),
    .B(n_10150_o_0),
    .C(n_10151_o_0),
    .Y(n_10511_o_0));
 AOI31xp33_ASAP7_75t_R n_10512 (.A1(n_10069_o_0),
    .A2(n_10085_o_0),
    .A3(n_10510_o_0),
    .B(n_10511_o_0),
    .Y(n_10512_o_0));
 AOI211xp5_ASAP7_75t_R n_10513 (.A1(n_10004_o_0),
    .A2(n_10509_o_0),
    .B(n_10512_o_0),
    .C(n_10146_o_0),
    .Y(n_10513_o_0));
 AOI31xp33_ASAP7_75t_R n_10514 (.A1(n_10077_o_0),
    .A2(n_10073_o_0),
    .A3(n_10225_o_0),
    .B(n_10359_o_0),
    .Y(n_10514_o_0));
 AOI321xp33_ASAP7_75t_R n_10515 (.A1(n_10214_o_0),
    .A2(n_10463_o_0),
    .A3(n_10004_o_0),
    .B1(n_10514_o_0),
    .B2(n_10150_o_0),
    .C(n_10067_o_0),
    .Y(n_10515_o_0));
 NOR3xp33_ASAP7_75t_R n_10516 (.A(n_10513_o_0),
    .B(n_10188_o_0),
    .C(n_10515_o_0),
    .Y(n_10516_o_0));
 AOI21xp33_ASAP7_75t_R n_10517 (.A1(n_10024_o_0),
    .A2(net61),
    .B(n_10160_o_0),
    .Y(n_10517_o_0));
 NOR3xp33_ASAP7_75t_R n_10518 (.A(n_10517_o_0),
    .B(n_10116_o_0),
    .C(n_10192_o_0),
    .Y(n_10518_o_0));
 OAI21xp33_ASAP7_75t_R n_10519 (.A1(n_10061_o_0),
    .A2(n_10178_o_0),
    .B(n_10067_o_0),
    .Y(n_10519_o_0));
 AOI21xp33_ASAP7_75t_R n_1052 (.A1(n_944_o_0),
    .A2(n_1051_o_0),
    .B(net16),
    .Y(n_1052_o_0));
 AOI21xp33_ASAP7_75t_R n_10520 (.A1(n_10085_o_0),
    .A2(n_10290_o_0),
    .B(n_10519_o_0),
    .Y(n_10520_o_0));
 OAI22xp33_ASAP7_75t_R n_10521 (.A1(n_10449_o_0),
    .A2(n_10200_o_0),
    .B1(n_10195_o_0),
    .B2(n_10242_o_0),
    .Y(n_10521_o_0));
 NOR3xp33_ASAP7_75t_R n_10522 (.A(n_10449_o_0),
    .B(n_10200_o_0),
    .C(n_10077_o_0),
    .Y(n_10522_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10523 (.A1(n_10521_o_0),
    .A2(n_10077_o_0),
    .B(n_10522_o_0),
    .C(n_10329_o_0),
    .Y(n_10523_o_0));
 OAI31xp33_ASAP7_75t_R n_10524 (.A1(n_10004_o_0),
    .A2(n_10518_o_0),
    .A3(n_10520_o_0),
    .B(n_10523_o_0),
    .Y(n_10524_o_0));
 AOI21xp33_ASAP7_75t_R n_10525 (.A1(net56),
    .A2(n_10087_o_0),
    .B(n_10085_o_0),
    .Y(n_10525_o_0));
 NOR2xp33_ASAP7_75t_R n_10526 (.A(n_10056_o_0),
    .B(n_10232_o_0),
    .Y(n_10526_o_0));
 AOI211xp5_ASAP7_75t_R n_10527 (.A1(n_10525_o_0),
    .A2(n_10319_o_0),
    .B(n_10526_o_0),
    .C(n_10308_o_0),
    .Y(n_10527_o_0));
 NOR3xp33_ASAP7_75t_R n_10528 (.A(n_10524_o_0),
    .B(n_10527_o_0),
    .C(n_10257_o_0),
    .Y(n_10528_o_0));
 INVx1_ASAP7_75t_R n_10529 (.A(n_10477_o_0),
    .Y(n_10529_o_0));
 OAI21xp33_ASAP7_75t_R n_1053 (.A1(n_877_o_0),
    .A2(n_1050_o_0),
    .B(n_1052_o_0),
    .Y(n_1053_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10530 (.A1(n_10213_o_0),
    .A2(n_10077_o_0),
    .B(n_10529_o_0),
    .C(n_10149_o_0),
    .Y(n_10530_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10531 (.A1(net24),
    .A2(net56),
    .B(n_10241_o_0),
    .C(n_10149_o_0),
    .Y(n_10531_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10532 (.A1(net24),
    .A2(n_10061_o_0),
    .B(n_10531_o_0),
    .C(n_10067_o_0),
    .Y(n_10532_o_0));
 AOI21xp33_ASAP7_75t_R n_10533 (.A1(n_10087_o_0),
    .A2(n_10203_o_0),
    .B(n_10005_o_0),
    .Y(n_10533_o_0));
 OAI21xp33_ASAP7_75t_R n_10534 (.A1(n_10170_o_0),
    .A2(n_10219_o_0),
    .B(n_10533_o_0),
    .Y(n_10534_o_0));
 OAI211xp5_ASAP7_75t_R n_10535 (.A1(n_10206_o_0),
    .A2(n_10489_o_0),
    .B(n_10268_o_0),
    .C(n_10150_o_0),
    .Y(n_10535_o_0));
 AOI21xp33_ASAP7_75t_R n_10536 (.A1(n_10534_o_0),
    .A2(n_10535_o_0),
    .B(n_10093_o_0),
    .Y(n_10536_o_0));
 AOI211xp5_ASAP7_75t_R n_10537 (.A1(n_10530_o_0),
    .A2(n_10532_o_0),
    .B(n_10536_o_0),
    .C(n_10313_o_0),
    .Y(n_10537_o_0));
 NOR2xp33_ASAP7_75t_R n_10538 (.A(n_10313_o_0),
    .B(n_9997_o_0),
    .Y(n_10538_o_0));
 OAI211xp5_ASAP7_75t_R n_10539 (.A1(n_10167_o_0),
    .A2(n_10129_o_0),
    .B(n_10005_o_0),
    .C(n_10208_o_0),
    .Y(n_10539_o_0));
 OAI211xp5_ASAP7_75t_R n_1054 (.A1(n_1049_o_0),
    .A2(net14),
    .B(n_903_o_0),
    .C(n_1053_o_0),
    .Y(n_1054_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10540 (.A1(n_10071_o_0),
    .A2(n_10125_o_0),
    .B(n_10466_o_0),
    .C(n_10539_o_0),
    .Y(n_10540_o_0));
 OAI21xp33_ASAP7_75t_R n_10541 (.A1(n_10245_o_0),
    .A2(n_10316_o_0),
    .B(n_10252_o_0),
    .Y(n_10541_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10542 (.A1(net56),
    .A2(n_10024_o_0),
    .B(net61),
    .C(n_10061_o_0),
    .Y(n_10542_o_0));
 AOI31xp33_ASAP7_75t_R n_10543 (.A1(n_10085_o_0),
    .A2(n_10380_o_0),
    .A3(n_10124_o_0),
    .B(n_10542_o_0),
    .Y(n_10543_o_0));
 AOI21xp33_ASAP7_75t_R n_10544 (.A1(n_10150_o_0),
    .A2(n_10543_o_0),
    .B(n_10067_o_0),
    .Y(n_10544_o_0));
 AOI21xp33_ASAP7_75t_R n_10545 (.A1(n_10541_o_0),
    .A2(n_10544_o_0),
    .B(n_10188_o_0),
    .Y(n_10545_o_0));
 OAI21xp33_ASAP7_75t_R n_10546 (.A1(n_10146_o_0),
    .A2(n_10540_o_0),
    .B(n_10545_o_0),
    .Y(n_10546_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10547 (.A1(n_10537_o_0),
    .A2(n_9997_o_0),
    .B(n_10538_o_0),
    .C(n_10546_o_0),
    .Y(n_10547_o_0));
 OAI31xp33_ASAP7_75t_R n_10548 (.A1(n_10102_o_0),
    .A2(n_10516_o_0),
    .A3(n_10528_o_0),
    .B(n_10547_o_0),
    .Y(n_10548_o_0));
 XOR2xp5_ASAP7_75t_R n_10549 (.A(_01009_),
    .B(_01096_),
    .Y(n_10549_o_0));
 AOI21xp33_ASAP7_75t_R n_1055 (.A1(n_886_o_0),
    .A2(n_908_o_0),
    .B(n_1041_o_0),
    .Y(n_1055_o_0));
 XNOR2xp5_ASAP7_75t_R n_10550 (.A(_01010_),
    .B(n_10549_o_0),
    .Y(n_10550_o_0));
 NOR2xp33_ASAP7_75t_R n_10551 (.A(n_3716_o_0),
    .B(n_10550_o_0),
    .Y(n_10551_o_0));
 NOR2xp33_ASAP7_75t_R n_10552 (.A(_00685_),
    .B(net),
    .Y(n_10552_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10553 (.A1(n_3716_o_0),
    .A2(n_10550_o_0),
    .B(n_10551_o_0),
    .C(net),
    .D(n_10552_o_0),
    .Y(n_10553_o_0));
 XNOR2xp5_ASAP7_75t_R n_10554 (.A(_00898_),
    .B(n_10553_o_0),
    .Y(n_10554_o_0));
 INVx1_ASAP7_75t_R n_10555 (.A(n_10554_o_0),
    .Y(n_10555_o_0));
 NOR2xp33_ASAP7_75t_R n_10556 (.A(n_3629_o_0),
    .B(n_8319_o_0),
    .Y(n_10556_o_0));
 XOR2xp5_ASAP7_75t_R n_10557 (.A(_01084_),
    .B(n_3643_o_0),
    .Y(n_10557_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10558 (.A1(n_3629_o_0),
    .A2(n_8319_o_0),
    .B(n_10556_o_0),
    .C(n_10557_o_0),
    .Y(n_10558_o_0));
 XNOR2xp5_ASAP7_75t_R n_10559 (.A(_01084_),
    .B(n_3643_o_0),
    .Y(n_10559_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1056 (.A1(net32),
    .A2(n_913_o_0),
    .B(n_1029_o_0),
    .C(n_877_o_0),
    .Y(n_1056_o_0));
 XNOR2xp5_ASAP7_75t_R n_10560 (.A(n_3629_o_0),
    .B(n_8323_o_0),
    .Y(n_10560_o_0));
 AOI21xp33_ASAP7_75t_R n_10561 (.A1(n_10559_o_0),
    .A2(n_10560_o_0),
    .B(n_3021_o_0),
    .Y(n_10561_o_0));
 AOI221xp5_ASAP7_75t_R n_10562 (.A1(n_3021_o_0),
    .A2(_00627_),
    .B1(n_10558_o_0),
    .B2(n_10561_o_0),
    .C(_00893_),
    .Y(n_10562_o_0));
 NAND2xp33_ASAP7_75t_R n_10563 (.A(_00627_),
    .B(net5),
    .Y(n_10563_o_0));
 OAI211xp5_ASAP7_75t_R n_10564 (.A1(n_10560_o_0),
    .A2(n_10559_o_0),
    .B(n_10561_o_0),
    .C(net),
    .Y(n_10564_o_0));
 INVx1_ASAP7_75t_R n_10565 (.A(_00893_),
    .Y(n_10565_o_0));
 AOI21xp33_ASAP7_75t_R n_10566 (.A1(n_10563_o_0),
    .A2(n_10564_o_0),
    .B(n_10565_o_0),
    .Y(n_10566_o_0));
 NOR2xp67_ASAP7_75t_R n_10567 (.A(n_10562_o_0),
    .B(n_10566_o_0),
    .Y(n_10567_o_0));
 INVx1_ASAP7_75t_R n_10568 (.A(_00894_),
    .Y(n_10568_o_0));
 XOR2xp5_ASAP7_75t_R n_10569 (.A(_01005_),
    .B(_01092_),
    .Y(n_10569_o_0));
 NOR3xp33_ASAP7_75t_R n_1057 (.A(n_934_o_0),
    .B(n_860_o_0),
    .C(n_878_o_0),
    .Y(n_1057_o_0));
 NAND2xp33_ASAP7_75t_R n_10570 (.A(_01085_),
    .B(n_10569_o_0),
    .Y(n_10570_o_0));
 OAI21xp33_ASAP7_75t_R n_10571 (.A1(_01085_),
    .A2(n_10569_o_0),
    .B(n_10570_o_0),
    .Y(n_10571_o_0));
 INVx1_ASAP7_75t_R n_10572 (.A(n_8306_o_0),
    .Y(n_10572_o_0));
 OAI211xp5_ASAP7_75t_R n_10573 (.A1(_01085_),
    .A2(n_10569_o_0),
    .B(n_10570_o_0),
    .C(n_10572_o_0),
    .Y(n_10573_o_0));
 INVx1_ASAP7_75t_R n_10574 (.A(n_10573_o_0),
    .Y(n_10574_o_0));
 NOR2xp33_ASAP7_75t_R n_10575 (.A(_00630_),
    .B(_00858_),
    .Y(n_10575_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10576 (.A1(n_8306_o_0),
    .A2(n_10571_o_0),
    .B(n_10574_o_0),
    .C(net77),
    .D(n_10575_o_0),
    .Y(n_10576_o_0));
 NAND2xp33_ASAP7_75t_R n_10577 (.A(n_8306_o_0),
    .B(n_10571_o_0),
    .Y(n_10577_o_0));
 INVx1_ASAP7_75t_R n_10578 (.A(n_10575_o_0),
    .Y(n_10578_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10579 (.A1(n_10573_o_0),
    .A2(n_10577_o_0),
    .B(n_3021_o_0),
    .C(n_10578_o_0),
    .D(n_10568_o_0),
    .Y(n_10579_o_0));
 OAI31xp33_ASAP7_75t_R n_1058 (.A1(n_903_o_0),
    .A2(n_1056_o_0),
    .A3(n_1057_o_0),
    .B(n_829_o_0),
    .Y(n_1058_o_0));
 AOI21x1_ASAP7_75t_R n_10580 (.A1(n_10568_o_0),
    .A2(n_10576_o_0),
    .B(n_10579_o_0),
    .Y(n_10580_o_0));
 XOR2xp5_ASAP7_75t_R n_10581 (.A(n_3667_o_0),
    .B(n_3643_o_0),
    .Y(n_10581_o_0));
 NOR2xp33_ASAP7_75t_R n_10582 (.A(_01098_),
    .B(n_10581_o_0),
    .Y(n_10582_o_0));
 NOR2xp33_ASAP7_75t_R n_10583 (.A(_00628_),
    .B(_00858_),
    .Y(n_10583_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10584 (.A1(n_10581_o_0),
    .A2(_01098_),
    .B(n_10582_o_0),
    .C(net39),
    .D(n_10583_o_0),
    .Y(n_10584_o_0));
 NAND2xp33_ASAP7_75t_R n_10585 (.A(n_3643_o_0),
    .B(n_3668_o_0),
    .Y(n_10585_o_0));
 INVx1_ASAP7_75t_R n_10586 (.A(_01098_),
    .Y(n_10586_o_0));
 OAI211xp5_ASAP7_75t_R n_10587 (.A1(n_3668_o_0),
    .A2(n_3643_o_0),
    .B(n_10585_o_0),
    .C(n_10586_o_0),
    .Y(n_10587_o_0));
 NAND2xp33_ASAP7_75t_R n_10588 (.A(_01098_),
    .B(n_10581_o_0),
    .Y(n_10588_o_0));
 INVx1_ASAP7_75t_R n_10589 (.A(n_10583_o_0),
    .Y(n_10589_o_0));
 AOI21xp33_ASAP7_75t_R n_1059 (.A1(n_1055_o_0),
    .A2(n_903_o_0),
    .B(n_1058_o_0),
    .Y(n_1059_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10590 (.A1(n_10587_o_0),
    .A2(n_10588_o_0),
    .B(net3),
    .C(n_10589_o_0),
    .D(_00892_),
    .Y(n_10590_o_0));
 AOI21x1_ASAP7_75t_R n_10591 (.A1(_00892_),
    .A2(n_10584_o_0),
    .B(n_10590_o_0),
    .Y(n_10591_o_0));
 NOR2xp33_ASAP7_75t_R n_10592 (.A(n_10580_o_0),
    .B(n_10591_o_0),
    .Y(n_10592_o_0));
 NAND2xp33_ASAP7_75t_R n_10593 (.A(n_10567_o_0),
    .B(n_10592_o_0),
    .Y(n_10593_o_0));
 OAI21xp33_ASAP7_75t_R n_10594 (.A1(n_10562_o_0),
    .A2(n_10566_o_0),
    .B(n_10591_o_0),
    .Y(n_10594_o_0));
 NAND2xp5_ASAP7_75t_R n_10595 (.A(n_10580_o_0),
    .B(n_10594_o_0),
    .Y(n_10595_o_0));
 INVx1_ASAP7_75t_R n_10596 (.A(_00895_),
    .Y(n_10596_o_0));
 XOR2xp5_ASAP7_75t_R n_10597 (.A(_01086_),
    .B(n_3614_o_0),
    .Y(n_10597_o_0));
 XNOR2xp5_ASAP7_75t_R n_10598 (.A(n_8298_o_0),
    .B(n_10597_o_0),
    .Y(n_10598_o_0));
 NOR2xp33_ASAP7_75t_R n_10599 (.A(_00688_),
    .B(_00858_),
    .Y(n_10599_o_0));
 INVx1_ASAP7_75t_R n_1060 (.A(n_956_o_0),
    .Y(n_1060_o_0));
 AOI21xp33_ASAP7_75t_R n_10600 (.A1(net77),
    .A2(n_10598_o_0),
    .B(n_10599_o_0),
    .Y(n_10600_o_0));
 XNOR2xp5_ASAP7_75t_R n_10601 (.A(n_8352_o_0),
    .B(n_10597_o_0),
    .Y(n_10601_o_0));
 INVx1_ASAP7_75t_R n_10602 (.A(n_10599_o_0),
    .Y(n_10602_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10603 (.A1(net1),
    .A2(n_10601_o_0),
    .B(n_10602_o_0),
    .C(n_10596_o_0),
    .Y(n_10603_o_0));
 AO21x1_ASAP7_75t_R n_10604 (.A1(n_10596_o_0),
    .A2(n_10600_o_0),
    .B(n_10603_o_0),
    .Y(n_10604_o_0));
 NAND3xp33_ASAP7_75t_R n_10605 (.A(n_10593_o_0),
    .B(n_10595_o_0),
    .C(n_10604_o_0),
    .Y(n_10605_o_0));
 XNOR2xp5_ASAP7_75t_R n_10606 (.A(_01087_),
    .B(n_3693_o_0),
    .Y(n_10606_o_0));
 NOR2xp33_ASAP7_75t_R n_10607 (.A(n_10606_o_0),
    .B(n_8375_o_0),
    .Y(n_10607_o_0));
 NOR2xp33_ASAP7_75t_R n_10608 (.A(_00687_),
    .B(net),
    .Y(n_10608_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10609 (.A1(n_8375_o_0),
    .A2(n_10606_o_0),
    .B(n_10607_o_0),
    .C(net),
    .D(n_10608_o_0),
    .Y(n_10609_o_0));
 NAND2xp33_ASAP7_75t_R n_1061 (.A(n_878_o_0),
    .B(n_903_o_0),
    .Y(n_1061_o_0));
 NAND2xp33_ASAP7_75t_R n_10610 (.A(_00896_),
    .B(n_10609_o_0),
    .Y(n_10610_o_0));
 OA21x2_ASAP7_75t_R n_10611 (.A1(_00896_),
    .A2(n_10609_o_0),
    .B(n_10610_o_0),
    .Y(n_10611_o_0));
 AOI22xp33_ASAP7_75t_R n_10612 (.A1(n_10561_o_0),
    .A2(n_10558_o_0),
    .B1(n_3021_o_0),
    .B2(_00627_),
    .Y(n_10612_o_0));
 INVx1_ASAP7_75t_R n_10613 (.A(n_10562_o_0),
    .Y(n_10613_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10614 (.A1(n_10612_o_0),
    .A2(n_10565_o_0),
    .B(n_10613_o_0),
    .C(n_10591_o_0),
    .Y(n_10614_o_0));
 INVx1_ASAP7_75t_R n_10615 (.A(n_10614_o_0),
    .Y(n_10615_o_0));
 NOR3xp33_ASAP7_75t_R n_10616 (.A(n_10615_o_0),
    .B(n_10604_o_0),
    .C(net43),
    .Y(n_10616_o_0));
 NOR2xp33_ASAP7_75t_R n_10617 (.A(n_10611_o_0),
    .B(n_10616_o_0),
    .Y(n_10617_o_0));
 INVx1_ASAP7_75t_R n_10618 (.A(n_10580_o_0),
    .Y(n_10618_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10619 (.A1(net1),
    .A2(n_10601_o_0),
    .B(n_10602_o_0),
    .C(_00895_),
    .Y(n_10619_o_0));
 OAI21xp33_ASAP7_75t_R n_1062 (.A1(n_881_o_0),
    .A2(n_918_o_0),
    .B(n_1051_o_0),
    .Y(n_1062_o_0));
 AO21x1_ASAP7_75t_R n_10620 (.A1(_00895_),
    .A2(n_10600_o_0),
    .B(n_10619_o_0),
    .Y(n_10620_o_0));
 OAI21xp33_ASAP7_75t_R n_10621 (.A1(n_10618_o_0),
    .A2(n_10594_o_0),
    .B(n_10620_o_0),
    .Y(n_10621_o_0));
 INVx1_ASAP7_75t_R n_10622 (.A(n_10621_o_0),
    .Y(n_10622_o_0));
 XNOR2xp5_ASAP7_75t_R n_10623 (.A(_00896_),
    .B(n_10609_o_0),
    .Y(n_10623_o_0));
 INVx1_ASAP7_75t_R n_10624 (.A(n_10623_o_0),
    .Y(n_10624_o_0));
 OAI31xp33_ASAP7_75t_R n_10625 (.A1(net43),
    .A2(n_10615_o_0),
    .A3(n_10620_o_0),
    .B(n_10624_o_0),
    .Y(n_10625_o_0));
 XNOR2xp5_ASAP7_75t_R n_10626 (.A(_01049_),
    .B(_01088_),
    .Y(n_10626_o_0));
 XNOR2xp5_ASAP7_75t_R n_10627 (.A(_01095_),
    .B(n_10626_o_0),
    .Y(n_10627_o_0));
 XOR2xp5_ASAP7_75t_R n_10628 (.A(_01008_),
    .B(_01009_),
    .Y(n_10628_o_0));
 NOR2xp33_ASAP7_75t_R n_10629 (.A(n_10628_o_0),
    .B(n_10627_o_0),
    .Y(n_10629_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1063 (.A1(n_1060_o_0),
    .A2(n_1061_o_0),
    .B(n_1062_o_0),
    .C(net16),
    .Y(n_1063_o_0));
 NOR2xp33_ASAP7_75t_R n_10630 (.A(_00686_),
    .B(net39),
    .Y(n_10630_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10631 (.A1(n_10627_o_0),
    .A2(n_10628_o_0),
    .B(n_10629_o_0),
    .C(net39),
    .D(n_10630_o_0),
    .Y(n_10631_o_0));
 XNOR2xp5_ASAP7_75t_R n_10632 (.A(_00897_),
    .B(n_10631_o_0),
    .Y(n_10632_o_0));
 INVx1_ASAP7_75t_R n_10633 (.A(n_10632_o_0),
    .Y(n_10633_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10634 (.A1(n_10622_o_0),
    .A2(n_10593_o_0),
    .B(n_10625_o_0),
    .C(n_10633_o_0),
    .Y(n_10634_o_0));
 AO21x1_ASAP7_75t_R n_10635 (.A1(n_10584_o_0),
    .A2(_00892_),
    .B(n_10590_o_0),
    .Y(n_10635_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10636 (.A1(n_10596_o_0),
    .A2(n_10600_o_0),
    .B(n_10603_o_0),
    .C(n_10580_o_0),
    .Y(n_10636_o_0));
 OAI211xp5_ASAP7_75t_R n_10637 (.A1(n_10591_o_0),
    .A2(n_10567_o_0),
    .B(n_10604_o_0),
    .C(n_10618_o_0),
    .Y(n_10637_o_0));
 OAI21xp33_ASAP7_75t_R n_10638 (.A1(n_10635_o_0),
    .A2(n_10636_o_0),
    .B(n_10637_o_0),
    .Y(n_10638_o_0));
 AOI21xp5_ASAP7_75t_R n_10639 (.A1(n_10596_o_0),
    .A2(n_10600_o_0),
    .B(n_10603_o_0),
    .Y(n_10639_o_0));
 NOR3xp33_ASAP7_75t_R n_1064 (.A(n_1059_o_0),
    .B(n_1063_o_0),
    .C(n_931_o_0),
    .Y(n_1064_o_0));
 NAND2xp33_ASAP7_75t_R n_10640 (.A(n_10580_o_0),
    .B(n_10639_o_0),
    .Y(n_10640_o_0));
 OAI21xp33_ASAP7_75t_R n_10641 (.A1(_00896_),
    .A2(n_10609_o_0),
    .B(n_10610_o_0),
    .Y(n_10641_o_0));
 OAI21xp33_ASAP7_75t_R n_10642 (.A1(n_10615_o_0),
    .A2(n_10640_o_0),
    .B(n_10641_o_0),
    .Y(n_10642_o_0));
 OAI21x1_ASAP7_75t_R n_10643 (.A1(n_10565_o_0),
    .A2(n_10612_o_0),
    .B(n_10613_o_0),
    .Y(n_10643_o_0));
 OAI21xp33_ASAP7_75t_R n_10644 (.A1(n_10591_o_0),
    .A2(n_10643_o_0),
    .B(n_10580_o_0),
    .Y(n_10644_o_0));
 OAI311xp33_ASAP7_75t_R n_10645 (.A1(n_10643_o_0),
    .A2(net43),
    .A3(n_10591_o_0),
    .B1(n_10620_o_0),
    .C1(n_10644_o_0),
    .Y(n_10645_o_0));
 INVx1_ASAP7_75t_R n_10646 (.A(n_10645_o_0),
    .Y(n_10646_o_0));
 NAND2xp33_ASAP7_75t_R n_10647 (.A(_00897_),
    .B(n_10631_o_0),
    .Y(n_10647_o_0));
 OAI21xp5_ASAP7_75t_R n_10648 (.A1(_00897_),
    .A2(n_10631_o_0),
    .B(n_10647_o_0),
    .Y(n_10648_o_0));
 NOR2xp33_ASAP7_75t_R n_10649 (.A(n_10580_o_0),
    .B(n_10643_o_0),
    .Y(n_10649_o_0));
 AOI311xp33_ASAP7_75t_R n_1065 (.A1(n_1048_o_0),
    .A2(n_1054_o_0),
    .A3(n_931_o_0),
    .B(n_972_o_0),
    .C(n_1064_o_0),
    .Y(n_1065_o_0));
 AOI21xp33_ASAP7_75t_R n_10650 (.A1(n_10587_o_0),
    .A2(n_10588_o_0),
    .B(net2),
    .Y(n_10650_o_0));
 INVx1_ASAP7_75t_R n_10651 (.A(_00892_),
    .Y(n_10651_o_0));
 AOI211xp5_ASAP7_75t_R n_10652 (.A1(n_10583_o_0),
    .A2(net2),
    .B(n_10650_o_0),
    .C(n_10651_o_0),
    .Y(n_10652_o_0));
 OAI22xp33_ASAP7_75t_R n_10653 (.A1(n_10652_o_0),
    .A2(n_10590_o_0),
    .B1(n_10566_o_0),
    .B2(n_10562_o_0),
    .Y(n_10653_o_0));
 OAI21xp5_ASAP7_75t_R n_10654 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(n_10653_o_0),
    .Y(n_10654_o_0));
 AOI21xp5_ASAP7_75t_R n_10655 (.A1(_00895_),
    .A2(n_10600_o_0),
    .B(n_10619_o_0),
    .Y(n_10655_o_0));
 OAI31xp33_ASAP7_75t_R n_10656 (.A1(net6),
    .A2(n_10654_o_0),
    .A3(n_10655_o_0),
    .B(n_10611_o_0),
    .Y(n_10656_o_0));
 AO21x1_ASAP7_75t_R n_10657 (.A1(n_10649_o_0),
    .A2(n_10604_o_0),
    .B(n_10656_o_0),
    .Y(n_10657_o_0));
 OAI311xp33_ASAP7_75t_R n_10658 (.A1(n_10638_o_0),
    .A2(n_10642_o_0),
    .A3(n_10646_o_0),
    .B1(n_10648_o_0),
    .C1(n_10657_o_0),
    .Y(n_10658_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10659 (.A1(n_10605_o_0),
    .A2(n_10617_o_0),
    .B(n_10634_o_0),
    .C(n_10658_o_0),
    .Y(n_10659_o_0));
 AO21x1_ASAP7_75t_R n_1066 (.A1(n_1040_o_0),
    .A2(n_972_o_0),
    .B(n_1065_o_0),
    .Y(n_1066_o_0));
 NOR2xp33_ASAP7_75t_R n_10660 (.A(n_10555_o_0),
    .B(n_10659_o_0),
    .Y(n_10660_o_0));
 NAND2xp33_ASAP7_75t_R n_10661 (.A(n_10635_o_0),
    .B(n_10567_o_0),
    .Y(n_10661_o_0));
 NOR2xp33_ASAP7_75t_R n_10662 (.A(n_10661_o_0),
    .B(n_10640_o_0),
    .Y(n_10662_o_0));
 NOR3xp33_ASAP7_75t_R n_10663 (.A(n_10643_o_0),
    .B(n_10635_o_0),
    .C(n_10580_o_0),
    .Y(n_10663_o_0));
 AOI211xp5_ASAP7_75t_R n_10664 (.A1(n_10568_o_0),
    .A2(n_10576_o_0),
    .B(n_10591_o_0),
    .C(n_10579_o_0),
    .Y(n_10664_o_0));
 NOR3xp33_ASAP7_75t_R n_10665 (.A(n_10663_o_0),
    .B(n_10664_o_0),
    .C(n_10639_o_0),
    .Y(n_10665_o_0));
 NOR3xp33_ASAP7_75t_R n_10666 (.A(n_10618_o_0),
    .B(n_10643_o_0),
    .C(n_10591_o_0),
    .Y(n_10666_o_0));
 INVx1_ASAP7_75t_R n_10667 (.A(n_10666_o_0),
    .Y(n_10667_o_0));
 AND2x2_ASAP7_75t_R n_10668 (.A(n_10568_o_0),
    .B(n_10576_o_0),
    .Y(n_10668_o_0));
 OAI211xp5_ASAP7_75t_R n_10669 (.A1(n_10668_o_0),
    .A2(n_10579_o_0),
    .B(n_10643_o_0),
    .C(n_10591_o_0),
    .Y(n_10669_o_0));
 INVx1_ASAP7_75t_R n_1067 (.A(n_890_o_0),
    .Y(n_1067_o_0));
 INVx1_ASAP7_75t_R n_10670 (.A(n_10636_o_0),
    .Y(n_10670_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10671 (.A1(n_10564_o_0),
    .A2(n_10563_o_0),
    .B(n_10565_o_0),
    .C(n_10613_o_0),
    .D(n_10591_o_0),
    .Y(n_10671_o_0));
 AOI211xp5_ASAP7_75t_R n_10672 (.A1(n_10591_o_0),
    .A2(n_10567_o_0),
    .B(n_10671_o_0),
    .C(n_10639_o_0),
    .Y(n_10672_o_0));
 AOI211xp5_ASAP7_75t_R n_10673 (.A1(n_10670_o_0),
    .A2(n_10654_o_0),
    .B(n_10672_o_0),
    .C(n_10641_o_0),
    .Y(n_10673_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10674 (.A1(n_10667_o_0),
    .A2(n_10669_o_0),
    .B(n_10604_o_0),
    .C(n_10673_o_0),
    .Y(n_10674_o_0));
 OAI31xp33_ASAP7_75t_R n_10675 (.A1(n_10611_o_0),
    .A2(n_10662_o_0),
    .A3(n_10665_o_0),
    .B(n_10674_o_0),
    .Y(n_10675_o_0));
 INVx1_ASAP7_75t_R n_10676 (.A(n_10592_o_0),
    .Y(n_10676_o_0));
 NOR2xp33_ASAP7_75t_R n_10677 (.A(n_10618_o_0),
    .B(n_10594_o_0),
    .Y(n_10677_o_0));
 NOR2xp33_ASAP7_75t_R n_10678 (.A(n_10639_o_0),
    .B(n_10677_o_0),
    .Y(n_10678_o_0));
 OAI211xp5_ASAP7_75t_R n_10679 (.A1(n_10643_o_0),
    .A2(n_10635_o_0),
    .B(n_10653_o_0),
    .C(n_10580_o_0),
    .Y(n_10679_o_0));
 AOI211xp5_ASAP7_75t_R n_1068 (.A1(n_860_o_0),
    .A2(net32),
    .B(n_877_o_0),
    .C(n_907_o_0),
    .Y(n_1068_o_0));
 AOI21xp33_ASAP7_75t_R n_10680 (.A1(n_10618_o_0),
    .A2(n_10567_o_0),
    .B(n_10655_o_0),
    .Y(n_10680_o_0));
 AOI21xp33_ASAP7_75t_R n_10681 (.A1(n_10679_o_0),
    .A2(n_10680_o_0),
    .B(n_10624_o_0),
    .Y(n_10681_o_0));
 INVx1_ASAP7_75t_R n_10682 (.A(n_10681_o_0),
    .Y(n_10682_o_0));
 NOR2xp33_ASAP7_75t_R n_10683 (.A(n_10591_o_0),
    .B(n_10643_o_0),
    .Y(n_10683_o_0));
 NOR2xp33_ASAP7_75t_R n_10684 (.A(n_10580_o_0),
    .B(n_10683_o_0),
    .Y(n_10684_o_0));
 AOI21xp33_ASAP7_75t_R n_10685 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(n_10618_o_0),
    .Y(n_10685_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10686 (.A1(net6),
    .A2(n_10614_o_0),
    .B(n_10685_o_0),
    .C(n_10639_o_0),
    .Y(n_10686_o_0));
 OAI211xp5_ASAP7_75t_R n_10687 (.A1(n_10684_o_0),
    .A2(n_10639_o_0),
    .B(n_10611_o_0),
    .C(n_10686_o_0),
    .Y(n_10687_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10688 (.A1(n_10676_o_0),
    .A2(n_10678_o_0),
    .B(n_10682_o_0),
    .C(n_10687_o_0),
    .Y(n_10688_o_0));
 AOI22xp33_ASAP7_75t_R n_10689 (.A1(n_10675_o_0),
    .A2(n_10648_o_0),
    .B1(n_10633_o_0),
    .B2(n_10688_o_0),
    .Y(n_10689_o_0));
 AOI21xp33_ASAP7_75t_R n_1069 (.A1(n_956_o_0),
    .A2(n_1067_o_0),
    .B(n_1068_o_0),
    .Y(n_1069_o_0));
 XOR2xp5_ASAP7_75t_R n_10690 (.A(_01010_),
    .B(_01097_),
    .Y(n_10690_o_0));
 XNOR2xp5_ASAP7_75t_R n_10691 (.A(_01011_),
    .B(n_10690_o_0),
    .Y(n_10691_o_0));
 NOR2xp33_ASAP7_75t_R n_10692 (.A(n_3607_o_0),
    .B(n_10691_o_0),
    .Y(n_10692_o_0));
 NOR2xp33_ASAP7_75t_R n_10693 (.A(_00684_),
    .B(net),
    .Y(n_10693_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10694 (.A1(n_3607_o_0),
    .A2(n_10691_o_0),
    .B(n_10692_o_0),
    .C(net),
    .D(n_10693_o_0),
    .Y(n_10694_o_0));
 NAND2xp33_ASAP7_75t_R n_10695 (.A(_00899_),
    .B(n_10694_o_0),
    .Y(n_10695_o_0));
 OAI21xp33_ASAP7_75t_R n_10696 (.A1(_00899_),
    .A2(n_10694_o_0),
    .B(n_10695_o_0),
    .Y(n_10696_o_0));
 INVx1_ASAP7_75t_R n_10697 (.A(n_10696_o_0),
    .Y(n_10697_o_0));
 OAI21xp33_ASAP7_75t_R n_10698 (.A1(n_10554_o_0),
    .A2(n_10689_o_0),
    .B(n_10697_o_0),
    .Y(n_10698_o_0));
 NAND2xp33_ASAP7_75t_R n_10699 (.A(_00898_),
    .B(n_10553_o_0),
    .Y(n_10699_o_0));
 AOI21xp33_ASAP7_75t_R n_1070 (.A1(n_1012_o_0),
    .A2(n_950_o_0),
    .B(n_954_o_0),
    .Y(n_1070_o_0));
 OAI21xp33_ASAP7_75t_R n_10700 (.A1(_00898_),
    .A2(n_10553_o_0),
    .B(n_10699_o_0),
    .Y(n_10700_o_0));
 INVx1_ASAP7_75t_R n_10701 (.A(n_10648_o_0),
    .Y(n_10701_o_0));
 NAND2xp33_ASAP7_75t_R n_10702 (.A(n_10580_o_0),
    .B(n_10635_o_0),
    .Y(n_10702_o_0));
 OAI21xp33_ASAP7_75t_R n_10703 (.A1(n_10643_o_0),
    .A2(n_10702_o_0),
    .B(n_10620_o_0),
    .Y(n_10703_o_0));
 OAI21xp33_ASAP7_75t_R n_10704 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(n_10618_o_0),
    .Y(n_10704_o_0));
 AOI31xp33_ASAP7_75t_R n_10705 (.A1(n_10604_o_0),
    .A2(n_10704_o_0),
    .A3(n_10702_o_0),
    .B(n_10641_o_0),
    .Y(n_10705_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10706 (.A1(net12),
    .A2(n_10643_o_0),
    .B(n_10703_o_0),
    .C(n_10705_o_0),
    .Y(n_10706_o_0));
 INVx1_ASAP7_75t_R n_10707 (.A(n_10706_o_0),
    .Y(n_10707_o_0));
 NOR2xp33_ASAP7_75t_R n_10708 (.A(n_10567_o_0),
    .B(n_10640_o_0),
    .Y(n_10708_o_0));
 NOR4xp25_ASAP7_75t_R n_10709 (.A(n_10665_o_0),
    .B(n_10708_o_0),
    .C(n_10611_o_0),
    .D(n_10616_o_0),
    .Y(n_10709_o_0));
 AOI21xp33_ASAP7_75t_R n_1071 (.A1(net15),
    .A2(n_1070_o_0),
    .B(n_903_o_0),
    .Y(n_1071_o_0));
 NAND3xp33_ASAP7_75t_R n_10710 (.A(n_10567_o_0),
    .B(n_10635_o_0),
    .C(n_10580_o_0),
    .Y(n_10710_o_0));
 INVx1_ASAP7_75t_R n_10711 (.A(n_10710_o_0),
    .Y(n_10711_o_0));
 NOR2xp33_ASAP7_75t_R n_10712 (.A(n_10655_o_0),
    .B(n_10664_o_0),
    .Y(n_10712_o_0));
 INVx1_ASAP7_75t_R n_10713 (.A(n_10712_o_0),
    .Y(n_10713_o_0));
 OAI31xp33_ASAP7_75t_R n_10714 (.A1(n_10639_o_0),
    .A2(n_10684_o_0),
    .A3(n_10711_o_0),
    .B(n_10713_o_0),
    .Y(n_10714_o_0));
 NAND3xp33_ASAP7_75t_R n_10715 (.A(n_10676_o_0),
    .B(n_10710_o_0),
    .C(n_10620_o_0),
    .Y(n_10715_o_0));
 INVx1_ASAP7_75t_R n_10716 (.A(n_10715_o_0),
    .Y(n_10716_o_0));
 AOI21xp33_ASAP7_75t_R n_10717 (.A1(n_10618_o_0),
    .A2(n_10654_o_0),
    .B(n_10639_o_0),
    .Y(n_10717_o_0));
 OAI21xp33_ASAP7_75t_R n_10718 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(n_10580_o_0),
    .Y(n_10718_o_0));
 AO21x1_ASAP7_75t_R n_10719 (.A1(n_10717_o_0),
    .A2(n_10718_o_0),
    .B(n_10641_o_0),
    .Y(n_10719_o_0));
 NOR2xp33_ASAP7_75t_R n_1072 (.A(n_989_o_0),
    .B(n_942_o_0),
    .Y(n_1072_o_0));
 OAI221xp5_ASAP7_75t_R n_10720 (.A1(n_10624_o_0),
    .A2(n_10714_o_0),
    .B1(n_10716_o_0),
    .B2(n_10719_o_0),
    .C(n_10633_o_0),
    .Y(n_10720_o_0));
 OAI31xp33_ASAP7_75t_R n_10721 (.A1(n_10701_o_0),
    .A2(n_10707_o_0),
    .A3(n_10709_o_0),
    .B(n_10720_o_0),
    .Y(n_10721_o_0));
 NAND2xp33_ASAP7_75t_R n_10722 (.A(n_10635_o_0),
    .B(n_10567_o_0),
    .Y(n_10722_o_0));
 NAND2xp33_ASAP7_75t_R n_10723 (.A(n_10580_o_0),
    .B(n_10591_o_0),
    .Y(n_10723_o_0));
 NAND3xp33_ASAP7_75t_R n_10724 (.A(n_10722_o_0),
    .B(n_10723_o_0),
    .C(n_10604_o_0),
    .Y(n_10724_o_0));
 NAND2xp33_ASAP7_75t_R n_10725 (.A(n_10635_o_0),
    .B(n_10643_o_0),
    .Y(n_10725_o_0));
 AOI21xp33_ASAP7_75t_R n_10726 (.A1(n_10618_o_0),
    .A2(n_10591_o_0),
    .B(n_10655_o_0),
    .Y(n_10726_o_0));
 NAND2xp33_ASAP7_75t_R n_10727 (.A(n_10725_o_0),
    .B(n_10726_o_0),
    .Y(n_10727_o_0));
 NAND4xp25_ASAP7_75t_R n_10728 (.A(n_10724_o_0),
    .B(n_10727_o_0),
    .C(n_10648_o_0),
    .D(n_10611_o_0),
    .Y(n_10728_o_0));
 OAI211xp5_ASAP7_75t_R n_10729 (.A1(n_10612_o_0),
    .A2(n_10565_o_0),
    .B(n_10591_o_0),
    .C(n_10613_o_0),
    .Y(n_10729_o_0));
 AOI31xp33_ASAP7_75t_R n_1073 (.A1(n_877_o_0),
    .A2(n_941_o_0),
    .A3(n_939_o_0),
    .B(n_1072_o_0),
    .Y(n_1073_o_0));
 NAND3xp33_ASAP7_75t_R n_10730 (.A(n_10620_o_0),
    .B(n_10729_o_0),
    .C(net43),
    .Y(n_10730_o_0));
 NAND3xp33_ASAP7_75t_R n_10731 (.A(n_10643_o_0),
    .B(n_10635_o_0),
    .C(n_10580_o_0),
    .Y(n_10731_o_0));
 OAI211xp5_ASAP7_75t_R n_10732 (.A1(n_10594_o_0),
    .A2(net43),
    .B(n_10731_o_0),
    .C(n_10604_o_0),
    .Y(n_10732_o_0));
 OAI311xp33_ASAP7_75t_R n_10733 (.A1(net43),
    .A2(n_10655_o_0),
    .A3(n_10654_o_0),
    .B1(n_10730_o_0),
    .C1(n_10732_o_0),
    .Y(n_10733_o_0));
 INVx1_ASAP7_75t_R n_10734 (.A(n_10725_o_0),
    .Y(n_10734_o_0));
 AOI211xp5_ASAP7_75t_R n_10735 (.A1(n_10598_o_0),
    .A2(net),
    .B(n_10596_o_0),
    .C(n_10599_o_0),
    .Y(n_10735_o_0));
 OAI22xp33_ASAP7_75t_R n_10736 (.A1(n_10635_o_0),
    .A2(n_10580_o_0),
    .B1(n_10619_o_0),
    .B2(n_10735_o_0),
    .Y(n_10736_o_0));
 OAI211xp5_ASAP7_75t_R n_10737 (.A1(n_10734_o_0),
    .A2(n_10736_o_0),
    .B(n_10724_o_0),
    .C(n_10611_o_0),
    .Y(n_10737_o_0));
 OAI31xp33_ASAP7_75t_R n_10738 (.A1(n_10648_o_0),
    .A2(n_10624_o_0),
    .A3(n_10733_o_0),
    .B(n_10737_o_0),
    .Y(n_10738_o_0));
 AOI21xp33_ASAP7_75t_R n_10739 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(n_10580_o_0),
    .Y(n_10739_o_0));
 AO21x1_ASAP7_75t_R n_1074 (.A1(n_881_o_0),
    .A2(n_935_o_0),
    .B(n_984_o_0),
    .Y(n_1074_o_0));
 INVx1_ASAP7_75t_R n_10740 (.A(n_10739_o_0),
    .Y(n_10740_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10741 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(n_10653_o_0),
    .C(n_10636_o_0),
    .Y(n_10741_o_0));
 AOI211xp5_ASAP7_75t_R n_10742 (.A1(n_10591_o_0),
    .A2(n_10643_o_0),
    .B(n_10655_o_0),
    .C(n_10618_o_0),
    .Y(n_10742_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10743 (.A1(n_10741_o_0),
    .A2(n_10672_o_0),
    .B(n_10731_o_0),
    .C(n_10742_o_0),
    .Y(n_10743_o_0));
 OAI21xp33_ASAP7_75t_R n_10744 (.A1(n_10740_o_0),
    .A2(n_10655_o_0),
    .B(n_10743_o_0),
    .Y(n_10744_o_0));
 AOI21xp33_ASAP7_75t_R n_10745 (.A1(net43),
    .A2(n_10654_o_0),
    .B(n_10620_o_0),
    .Y(n_10745_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10746 (.A1(n_10591_o_0),
    .A2(n_10567_o_0),
    .B(n_10671_o_0),
    .C(n_10618_o_0),
    .Y(n_10746_o_0));
 AOI31xp33_ASAP7_75t_R n_10747 (.A1(n_10643_o_0),
    .A2(n_10639_o_0),
    .A3(net43),
    .B(n_10623_o_0),
    .Y(n_10747_o_0));
 OAI21xp33_ASAP7_75t_R n_10748 (.A1(n_10604_o_0),
    .A2(n_10746_o_0),
    .B(n_10747_o_0),
    .Y(n_10748_o_0));
 OAI21xp33_ASAP7_75t_R n_10749 (.A1(n_10745_o_0),
    .A2(n_10748_o_0),
    .B(n_10632_o_0),
    .Y(n_10749_o_0));
 OAI221xp5_ASAP7_75t_R n_1075 (.A1(n_989_o_0),
    .A2(n_991_o_0),
    .B1(n_877_o_0),
    .B2(n_1074_o_0),
    .C(n_891_o_0),
    .Y(n_1075_o_0));
 AOI21xp33_ASAP7_75t_R n_10750 (.A1(n_10641_o_0),
    .A2(n_10744_o_0),
    .B(n_10749_o_0),
    .Y(n_10750_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10751 (.A1(n_10728_o_0),
    .A2(n_10738_o_0),
    .B(n_10750_o_0),
    .C(n_10554_o_0),
    .D(n_10697_o_0),
    .Y(n_10751_o_0));
 OAI21xp33_ASAP7_75t_R n_10752 (.A1(n_10700_o_0),
    .A2(n_10721_o_0),
    .B(n_10751_o_0),
    .Y(n_10752_o_0));
 OAI21xp33_ASAP7_75t_R n_10753 (.A1(n_10660_o_0),
    .A2(n_10698_o_0),
    .B(n_10752_o_0),
    .Y(n_10753_o_0));
 XNOR2xp5_ASAP7_75t_R n_10754 (.A(_00899_),
    .B(n_10694_o_0),
    .Y(n_10754_o_0));
 AOI21xp33_ASAP7_75t_R n_10755 (.A1(net43),
    .A2(n_10654_o_0),
    .B(n_10736_o_0),
    .Y(n_10755_o_0));
 AOI31xp33_ASAP7_75t_R n_10756 (.A1(n_10604_o_0),
    .A2(n_10676_o_0),
    .A3(n_10729_o_0),
    .B(n_10755_o_0),
    .Y(n_10756_o_0));
 OAI21xp33_ASAP7_75t_R n_10757 (.A1(n_10619_o_0),
    .A2(n_10735_o_0),
    .B(n_10723_o_0),
    .Y(n_10757_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10758 (.A1(net12),
    .A2(n_10615_o_0),
    .B(n_10757_o_0),
    .C(n_10611_o_0),
    .Y(n_10758_o_0));
 AOI21xp33_ASAP7_75t_R n_10759 (.A1(n_10667_o_0),
    .A2(n_10717_o_0),
    .B(n_10758_o_0),
    .Y(n_10759_o_0));
 OAI21xp33_ASAP7_75t_R n_1076 (.A1(n_1073_o_0),
    .A2(net14),
    .B(n_1075_o_0),
    .Y(n_1076_o_0));
 AOI21xp33_ASAP7_75t_R n_10760 (.A1(n_10623_o_0),
    .A2(n_10756_o_0),
    .B(n_10759_o_0),
    .Y(n_10760_o_0));
 NAND2xp33_ASAP7_75t_R n_10761 (.A(n_10580_o_0),
    .B(n_10567_o_0),
    .Y(n_10761_o_0));
 AOI21xp33_ASAP7_75t_R n_10762 (.A1(n_10604_o_0),
    .A2(n_10761_o_0),
    .B(n_10641_o_0),
    .Y(n_10762_o_0));
 INVx1_ASAP7_75t_R n_10763 (.A(n_10762_o_0),
    .Y(n_10763_o_0));
 NAND2xp33_ASAP7_75t_R n_10764 (.A(n_10643_o_0),
    .B(n_10618_o_0),
    .Y(n_10764_o_0));
 OAI21xp33_ASAP7_75t_R n_10765 (.A1(n_10661_o_0),
    .A2(n_10640_o_0),
    .B(n_10764_o_0),
    .Y(n_10765_o_0));
 OAI211xp5_ASAP7_75t_R n_10766 (.A1(n_10612_o_0),
    .A2(n_10565_o_0),
    .B(n_10591_o_0),
    .C(n_10613_o_0),
    .Y(n_10766_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10767 (.A1(n_10766_o_0),
    .A2(n_10653_o_0),
    .B(n_10618_o_0),
    .C(n_10604_o_0),
    .Y(n_10767_o_0));
 INVx1_ASAP7_75t_R n_10768 (.A(n_10704_o_0),
    .Y(n_10768_o_0));
 OAI211xp5_ASAP7_75t_R n_10769 (.A1(n_10767_o_0),
    .A2(n_10768_o_0),
    .B(n_10645_o_0),
    .C(n_10623_o_0),
    .Y(n_10769_o_0));
 AO21x1_ASAP7_75t_R n_1077 (.A1(n_1076_o_0),
    .A2(n_903_o_0),
    .B(n_931_o_0),
    .Y(n_1077_o_0));
 OAI211xp5_ASAP7_75t_R n_10770 (.A1(n_10763_o_0),
    .A2(n_10765_o_0),
    .B(n_10769_o_0),
    .C(n_10700_o_0),
    .Y(n_10770_o_0));
 OAI21xp33_ASAP7_75t_R n_10771 (.A1(n_10554_o_0),
    .A2(n_10760_o_0),
    .B(n_10770_o_0),
    .Y(n_10771_o_0));
 INVx1_ASAP7_75t_R n_10772 (.A(n_10684_o_0),
    .Y(n_10772_o_0));
 AOI211xp5_ASAP7_75t_R n_10773 (.A1(n_10654_o_0),
    .A2(net6),
    .B(n_10639_o_0),
    .C(n_10664_o_0),
    .Y(n_10773_o_0));
 AOI31xp33_ASAP7_75t_R n_10774 (.A1(n_10620_o_0),
    .A2(n_10772_o_0),
    .A3(n_10723_o_0),
    .B(n_10773_o_0),
    .Y(n_10774_o_0));
 AO21x1_ASAP7_75t_R n_10775 (.A1(n_10680_o_0),
    .A2(n_10725_o_0),
    .B(n_10624_o_0),
    .Y(n_10775_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10776 (.A1(n_10722_o_0),
    .A2(n_10670_o_0),
    .B(n_10775_o_0),
    .C(n_10700_o_0),
    .Y(n_10776_o_0));
 OAI21xp33_ASAP7_75t_R n_10777 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(n_10618_o_0),
    .Y(n_10777_o_0));
 INVx1_ASAP7_75t_R n_10778 (.A(n_10777_o_0),
    .Y(n_10778_o_0));
 AOI211xp5_ASAP7_75t_R n_10779 (.A1(n_10580_o_0),
    .A2(n_10635_o_0),
    .B(n_10639_o_0),
    .C(n_10643_o_0),
    .Y(n_10779_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1078 (.A1(net15),
    .A2(n_1069_o_0),
    .B(n_1071_o_0),
    .C(n_1077_o_0),
    .Y(n_1078_o_0));
 AO21x1_ASAP7_75t_R n_10780 (.A1(n_10620_o_0),
    .A2(n_10778_o_0),
    .B(n_10779_o_0),
    .Y(n_10780_o_0));
 OAI211xp5_ASAP7_75t_R n_10781 (.A1(n_10643_o_0),
    .A2(n_10635_o_0),
    .B(n_10618_o_0),
    .C(n_10653_o_0),
    .Y(n_10781_o_0));
 AOI31xp33_ASAP7_75t_R n_10782 (.A1(n_10591_o_0),
    .A2(n_10580_o_0),
    .A3(n_10567_o_0),
    .B(n_10639_o_0),
    .Y(n_10782_o_0));
 AOI21xp33_ASAP7_75t_R n_10783 (.A1(n_10781_o_0),
    .A2(n_10782_o_0),
    .B(n_10624_o_0),
    .Y(n_10783_o_0));
 OAI31xp33_ASAP7_75t_R n_10784 (.A1(n_10604_o_0),
    .A2(n_10661_o_0),
    .A3(net43),
    .B(n_10783_o_0),
    .Y(n_10784_o_0));
 OAI211xp5_ASAP7_75t_R n_10785 (.A1(n_10641_o_0),
    .A2(n_10780_o_0),
    .B(n_10784_o_0),
    .C(n_10555_o_0),
    .Y(n_10785_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10786 (.A1(n_10774_o_0),
    .A2(n_10611_o_0),
    .B(n_10776_o_0),
    .C(n_10785_o_0),
    .Y(n_10786_o_0));
 OAI22xp33_ASAP7_75t_R n_10787 (.A1(n_10771_o_0),
    .A2(n_10633_o_0),
    .B1(n_10648_o_0),
    .B2(n_10786_o_0),
    .Y(n_10787_o_0));
 OAI21xp33_ASAP7_75t_R n_10788 (.A1(n_10567_o_0),
    .A2(n_10618_o_0),
    .B(n_10604_o_0),
    .Y(n_10788_o_0));
 OAI21xp33_ASAP7_75t_R n_10789 (.A1(n_10788_o_0),
    .A2(n_10684_o_0),
    .B(n_10701_o_0),
    .Y(n_10789_o_0));
 OAI31xp33_ASAP7_75t_R n_1079 (.A1(n_878_o_0),
    .A2(n_907_o_0),
    .A3(n_913_o_0),
    .B(n_829_o_0),
    .Y(n_1079_o_0));
 AOI21xp33_ASAP7_75t_R n_10790 (.A1(n_10653_o_0),
    .A2(n_10766_o_0),
    .B(n_10580_o_0),
    .Y(n_10790_o_0));
 NOR2xp33_ASAP7_75t_R n_10791 (.A(n_10580_o_0),
    .B(n_10635_o_0),
    .Y(n_10791_o_0));
 INVx1_ASAP7_75t_R n_10792 (.A(n_10791_o_0),
    .Y(n_10792_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10793 (.A1(n_10643_o_0),
    .A2(n_10792_o_0),
    .B(n_10712_o_0),
    .C(n_10633_o_0),
    .Y(n_10793_o_0));
 OAI21xp33_ASAP7_75t_R n_10794 (.A1(n_10639_o_0),
    .A2(n_10790_o_0),
    .B(n_10793_o_0),
    .Y(n_10794_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10795 (.A1(n_10731_o_0),
    .A2(n_10726_o_0),
    .B(n_10789_o_0),
    .C(n_10794_o_0),
    .Y(n_10795_o_0));
 INVx1_ASAP7_75t_R n_10796 (.A(n_10700_o_0),
    .Y(n_10796_o_0));
 NAND2xp33_ASAP7_75t_R n_10797 (.A(net43),
    .B(n_10643_o_0),
    .Y(n_10797_o_0));
 NOR2xp33_ASAP7_75t_R n_10798 (.A(n_10663_o_0),
    .B(n_10621_o_0),
    .Y(n_10798_o_0));
 AOI31xp33_ASAP7_75t_R n_10799 (.A1(n_10648_o_0),
    .A2(n_10604_o_0),
    .A3(n_10797_o_0),
    .B(n_10798_o_0),
    .Y(n_10799_o_0));
 NOR3xp33_ASAP7_75t_R n_1080 (.A(n_1060_o_0),
    .B(n_877_o_0),
    .C(n_982_o_0),
    .Y(n_1080_o_0));
 OAI22xp33_ASAP7_75t_R n_10800 (.A1(n_10795_o_0),
    .A2(n_10554_o_0),
    .B1(n_10796_o_0),
    .B2(n_10799_o_0),
    .Y(n_10800_o_0));
 OAI211xp5_ASAP7_75t_R n_10801 (.A1(n_10580_o_0),
    .A2(n_10635_o_0),
    .B(n_10604_o_0),
    .C(n_10567_o_0),
    .Y(n_10801_o_0));
 NAND2xp33_ASAP7_75t_R n_10802 (.A(n_10632_o_0),
    .B(n_10801_o_0),
    .Y(n_10802_o_0));
 NOR2xp33_ASAP7_75t_R n_10803 (.A(n_10655_o_0),
    .B(n_10592_o_0),
    .Y(n_10803_o_0));
 INVx1_ASAP7_75t_R n_10804 (.A(n_10803_o_0),
    .Y(n_10804_o_0));
 AOI21xp33_ASAP7_75t_R n_10805 (.A1(n_10591_o_0),
    .A2(n_10567_o_0),
    .B(net43),
    .Y(n_10805_o_0));
 AOI21xp33_ASAP7_75t_R n_10806 (.A1(n_10567_o_0),
    .A2(n_10635_o_0),
    .B(n_10618_o_0),
    .Y(n_10806_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10807 (.A1(n_10805_o_0),
    .A2(n_10806_o_0),
    .B(n_10604_o_0),
    .C(n_10648_o_0),
    .Y(n_10807_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10808 (.A1(net43),
    .A2(n_10614_o_0),
    .B(n_10804_o_0),
    .C(n_10807_o_0),
    .D(n_10796_o_0),
    .Y(n_10808_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10809 (.A1(n_10726_o_0),
    .A2(n_10761_o_0),
    .B(n_10802_o_0),
    .C(n_10808_o_0),
    .Y(n_10809_o_0));
 NAND3xp33_ASAP7_75t_R n_1081 (.A(n_882_o_0),
    .B(n_990_o_0),
    .C(n_878_o_0),
    .Y(n_1081_o_0));
 AOI31xp33_ASAP7_75t_R n_10810 (.A1(n_10766_o_0),
    .A2(net43),
    .A3(n_10653_o_0),
    .B(n_10620_o_0),
    .Y(n_10810_o_0));
 AOI21xp33_ASAP7_75t_R n_10811 (.A1(n_10591_o_0),
    .A2(n_10580_o_0),
    .B(n_10604_o_0),
    .Y(n_10811_o_0));
 NAND2xp33_ASAP7_75t_R n_10812 (.A(n_10618_o_0),
    .B(n_10620_o_0),
    .Y(n_10812_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10813 (.A1(n_10637_o_0),
    .A2(n_10810_o_0),
    .B(n_10811_o_0),
    .C(n_10812_o_0),
    .D(n_10615_o_0),
    .Y(n_10813_o_0));
 AOI211xp5_ASAP7_75t_R n_10814 (.A1(n_10810_o_0),
    .A2(n_10637_o_0),
    .B(n_10614_o_0),
    .C(n_10811_o_0),
    .Y(n_10814_o_0));
 INVx1_ASAP7_75t_R n_10815 (.A(n_10654_o_0),
    .Y(n_10815_o_0));
 OAI21xp33_ASAP7_75t_R n_10816 (.A1(n_10618_o_0),
    .A2(n_10729_o_0),
    .B(n_10604_o_0),
    .Y(n_10816_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10817 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(n_10618_o_0),
    .C(n_10655_o_0),
    .Y(n_10817_o_0));
 INVx1_ASAP7_75t_R n_10818 (.A(n_10685_o_0),
    .Y(n_10818_o_0));
 AOI21xp33_ASAP7_75t_R n_10819 (.A1(n_10817_o_0),
    .A2(n_10818_o_0),
    .B(n_10633_o_0),
    .Y(n_10819_o_0));
 OAI31xp33_ASAP7_75t_R n_1082 (.A1(n_878_o_0),
    .A2(n_934_o_0),
    .A3(n_1006_o_0),
    .B(n_1081_o_0),
    .Y(n_1082_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10820 (.A1(net6),
    .A2(n_10815_o_0),
    .B(n_10816_o_0),
    .C(n_10819_o_0),
    .D(n_10554_o_0),
    .Y(n_10820_o_0));
 OAI31xp33_ASAP7_75t_R n_10821 (.A1(n_10648_o_0),
    .A2(n_10813_o_0),
    .A3(n_10814_o_0),
    .B(n_10820_o_0),
    .Y(n_10821_o_0));
 AOI31xp33_ASAP7_75t_R n_10822 (.A1(n_10611_o_0),
    .A2(n_10809_o_0),
    .A3(n_10821_o_0),
    .B(n_10697_o_0),
    .Y(n_10822_o_0));
 OAI21xp33_ASAP7_75t_R n_10823 (.A1(n_10624_o_0),
    .A2(n_10800_o_0),
    .B(n_10822_o_0),
    .Y(n_10823_o_0));
 OAI21xp33_ASAP7_75t_R n_10824 (.A1(n_10754_o_0),
    .A2(n_10787_o_0),
    .B(n_10823_o_0),
    .Y(n_10824_o_0));
 INVx1_ASAP7_75t_R n_10825 (.A(n_10594_o_0),
    .Y(n_10825_o_0));
 AOI211xp5_ASAP7_75t_R n_10826 (.A1(n_10591_o_0),
    .A2(n_10580_o_0),
    .B(n_10639_o_0),
    .C(n_10643_o_0),
    .Y(n_10826_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10827 (.A1(net12),
    .A2(n_10825_o_0),
    .B(n_10666_o_0),
    .C(n_10639_o_0),
    .D(n_10826_o_0),
    .Y(n_10827_o_0));
 OAI311xp33_ASAP7_75t_R n_10828 (.A1(n_10635_o_0),
    .A2(n_10618_o_0),
    .A3(n_10643_o_0),
    .B1(n_10620_o_0),
    .C1(n_10669_o_0),
    .Y(n_10828_o_0));
 OAI31xp33_ASAP7_75t_R n_10829 (.A1(n_10639_o_0),
    .A2(n_10791_o_0),
    .A3(n_10666_o_0),
    .B(n_10828_o_0),
    .Y(n_10829_o_0));
 AOI21xp33_ASAP7_75t_R n_1083 (.A1(net15),
    .A2(n_1082_o_0),
    .B(n_903_o_0),
    .Y(n_1083_o_0));
 AO22x1_ASAP7_75t_R n_10830 (.A1(n_10641_o_0),
    .A2(n_10827_o_0),
    .B1(n_10829_o_0),
    .B2(n_10624_o_0),
    .Y(n_10830_o_0));
 AO22x1_ASAP7_75t_R n_10831 (.A1(n_10595_o_0),
    .A2(n_10803_o_0),
    .B1(n_10717_o_0),
    .B2(n_10679_o_0),
    .Y(n_10831_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10832 (.A1(net43),
    .A2(n_10643_o_0),
    .B(n_10635_o_0),
    .C(n_10620_o_0),
    .D(n_10641_o_0),
    .Y(n_10832_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10833 (.A1(n_10825_o_0),
    .A2(net12),
    .B(n_10788_o_0),
    .C(n_10832_o_0),
    .Y(n_10833_o_0));
 NAND2xp33_ASAP7_75t_R n_10834 (.A(n_10633_o_0),
    .B(n_10833_o_0),
    .Y(n_10834_o_0));
 AOI21xp33_ASAP7_75t_R n_10835 (.A1(n_10623_o_0),
    .A2(n_10831_o_0),
    .B(n_10834_o_0),
    .Y(n_10835_o_0));
 AOI21xp33_ASAP7_75t_R n_10836 (.A1(n_10648_o_0),
    .A2(n_10830_o_0),
    .B(n_10835_o_0),
    .Y(n_10836_o_0));
 INVx1_ASAP7_75t_R n_10837 (.A(n_10754_o_0),
    .Y(n_10837_o_0));
 NOR3xp33_ASAP7_75t_R n_10838 (.A(n_10643_o_0),
    .B(n_10580_o_0),
    .C(n_10591_o_0),
    .Y(n_10838_o_0));
 OAI21xp33_ASAP7_75t_R n_10839 (.A1(n_10838_o_0),
    .A2(n_10767_o_0),
    .B(n_10623_o_0),
    .Y(n_10839_o_0));
 OAI21xp33_ASAP7_75t_R n_1084 (.A1(n_1079_o_0),
    .A2(n_1080_o_0),
    .B(n_1083_o_0),
    .Y(n_1084_o_0));
 AOI21xp33_ASAP7_75t_R n_10840 (.A1(n_10649_o_0),
    .A2(n_10620_o_0),
    .B(n_10839_o_0),
    .Y(n_10840_o_0));
 OAI21xp33_ASAP7_75t_R n_10841 (.A1(n_10592_o_0),
    .A2(n_10788_o_0),
    .B(n_10611_o_0),
    .Y(n_10841_o_0));
 AOI21xp33_ASAP7_75t_R n_10842 (.A1(n_10679_o_0),
    .A2(n_10680_o_0),
    .B(n_10841_o_0),
    .Y(n_10842_o_0));
 NAND2xp33_ASAP7_75t_R n_10843 (.A(n_10618_o_0),
    .B(n_10594_o_0),
    .Y(n_10843_o_0));
 AOI211xp5_ASAP7_75t_R n_10844 (.A1(n_10591_o_0),
    .A2(n_10580_o_0),
    .B(n_10655_o_0),
    .C(n_10567_o_0),
    .Y(n_10844_o_0));
 AOI31xp33_ASAP7_75t_R n_10845 (.A1(n_10604_o_0),
    .A2(n_10679_o_0),
    .A3(n_10843_o_0),
    .B(n_10844_o_0),
    .Y(n_10845_o_0));
 NAND3xp33_ASAP7_75t_R n_10846 (.A(n_10845_o_0),
    .B(n_10624_o_0),
    .C(n_10648_o_0),
    .Y(n_10846_o_0));
 OAI211xp5_ASAP7_75t_R n_10847 (.A1(n_10643_o_0),
    .A2(n_10580_o_0),
    .B(n_10725_o_0),
    .C(n_10604_o_0),
    .Y(n_10847_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10848 (.A1(net43),
    .A2(n_10643_o_0),
    .B(n_10655_o_0),
    .C(n_10847_o_0),
    .Y(n_10848_o_0));
 NAND3xp33_ASAP7_75t_R n_10849 (.A(n_10848_o_0),
    .B(n_10648_o_0),
    .C(n_10623_o_0),
    .Y(n_10849_o_0));
 INVx1_ASAP7_75t_R n_1085 (.A(n_982_o_0),
    .Y(n_1085_o_0));
 OAI311xp33_ASAP7_75t_R n_10850 (.A1(n_10632_o_0),
    .A2(n_10840_o_0),
    .A3(n_10842_o_0),
    .B1(n_10846_o_0),
    .C1(n_10849_o_0),
    .Y(n_10850_o_0));
 OAI22xp33_ASAP7_75t_R n_10851 (.A1(n_10836_o_0),
    .A2(n_10837_o_0),
    .B1(n_10696_o_0),
    .B2(n_10850_o_0),
    .Y(n_10851_o_0));
 NAND2xp33_ASAP7_75t_R n_10852 (.A(n_10580_o_0),
    .B(n_10643_o_0),
    .Y(n_10852_o_0));
 AOI211xp5_ASAP7_75t_R n_10853 (.A1(net43),
    .A2(n_10614_o_0),
    .B(n_10791_o_0),
    .C(n_10639_o_0),
    .Y(n_10853_o_0));
 AOI31xp33_ASAP7_75t_R n_10854 (.A1(n_10620_o_0),
    .A2(n_10781_o_0),
    .A3(n_10852_o_0),
    .B(n_10853_o_0),
    .Y(n_10854_o_0));
 NOR2xp33_ASAP7_75t_R n_10855 (.A(n_10632_o_0),
    .B(n_10623_o_0),
    .Y(n_10855_o_0));
 INVx1_ASAP7_75t_R n_10856 (.A(n_10855_o_0),
    .Y(n_10856_o_0));
 AOI21xp33_ASAP7_75t_R n_10857 (.A1(n_10618_o_0),
    .A2(n_10661_o_0),
    .B(n_10604_o_0),
    .Y(n_10857_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10858 (.A1(n_10635_o_0),
    .A2(n_10618_o_0),
    .B(n_10567_o_0),
    .C(n_10639_o_0),
    .Y(n_10858_o_0));
 AOI21xp33_ASAP7_75t_R n_10859 (.A1(n_10718_o_0),
    .A2(n_10857_o_0),
    .B(n_10858_o_0),
    .Y(n_10859_o_0));
 OAI211xp5_ASAP7_75t_R n_1086 (.A1(n_957_o_0),
    .A2(n_881_o_0),
    .B(n_877_o_0),
    .C(n_1085_o_0),
    .Y(n_1086_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10860 (.A1(n_10661_o_0),
    .A2(net43),
    .B(n_10838_o_0),
    .C(n_10655_o_0),
    .Y(n_10860_o_0));
 AOI21xp33_ASAP7_75t_R n_10861 (.A1(n_10681_o_0),
    .A2(n_10860_o_0),
    .B(n_10701_o_0),
    .Y(n_10861_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10862 (.A1(n_10664_o_0),
    .A2(n_10567_o_0),
    .B(n_10655_o_0),
    .C(n_10623_o_0),
    .Y(n_10862_o_0));
 AOI211xp5_ASAP7_75t_R n_10863 (.A1(n_10704_o_0),
    .A2(n_10782_o_0),
    .B(n_10862_o_0),
    .C(n_10648_o_0),
    .Y(n_10863_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10864 (.A1(n_10623_o_0),
    .A2(n_10859_o_0),
    .B(n_10861_o_0),
    .C(n_10863_o_0),
    .Y(n_10864_o_0));
 OAI21xp33_ASAP7_75t_R n_10865 (.A1(n_10854_o_0),
    .A2(n_10856_o_0),
    .B(n_10864_o_0),
    .Y(n_10865_o_0));
 OA21x2_ASAP7_75t_R n_10866 (.A1(n_10639_o_0),
    .A2(n_10649_o_0),
    .B(n_10703_o_0),
    .Y(n_10866_o_0));
 OAI31xp33_ASAP7_75t_R n_10867 (.A1(n_10618_o_0),
    .A2(n_10604_o_0),
    .A3(n_10643_o_0),
    .B(n_10624_o_0),
    .Y(n_10867_o_0));
 OAI21xp33_ASAP7_75t_R n_10868 (.A1(n_10858_o_0),
    .A2(n_10867_o_0),
    .B(n_10648_o_0),
    .Y(n_10868_o_0));
 AOI21xp33_ASAP7_75t_R n_10869 (.A1(n_10623_o_0),
    .A2(n_10866_o_0),
    .B(n_10868_o_0),
    .Y(n_10869_o_0));
 OAI31xp33_ASAP7_75t_R n_1087 (.A1(n_907_o_0),
    .A2(n_984_o_0),
    .A3(n_877_o_0),
    .B(n_1086_o_0),
    .Y(n_1087_o_0));
 NOR2xp33_ASAP7_75t_R n_10870 (.A(n_10580_o_0),
    .B(n_10635_o_0),
    .Y(n_10870_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10871 (.A1(n_10643_o_0),
    .A2(n_10792_o_0),
    .B(n_10622_o_0),
    .C(n_10641_o_0),
    .Y(n_10871_o_0));
 OAI31xp33_ASAP7_75t_R n_10872 (.A1(net43),
    .A2(n_10614_o_0),
    .A3(n_10655_o_0),
    .B(n_10623_o_0),
    .Y(n_10872_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10873 (.A1(n_10717_o_0),
    .A2(n_10644_o_0),
    .B(n_10872_o_0),
    .C(n_10633_o_0),
    .Y(n_10873_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10874 (.A1(n_10816_o_0),
    .A2(n_10870_o_0),
    .B(n_10871_o_0),
    .C(n_10873_o_0),
    .Y(n_10874_o_0));
 OAI31xp33_ASAP7_75t_R n_10875 (.A1(n_10869_o_0),
    .A2(n_10874_o_0),
    .A3(n_10696_o_0),
    .B(n_10700_o_0),
    .Y(n_10875_o_0));
 AO21x1_ASAP7_75t_R n_10876 (.A1(n_10865_o_0),
    .A2(n_10754_o_0),
    .B(n_10875_o_0),
    .Y(n_10876_o_0));
 OAI21xp33_ASAP7_75t_R n_10877 (.A1(n_10554_o_0),
    .A2(n_10851_o_0),
    .B(n_10876_o_0),
    .Y(n_10877_o_0));
 AOI21xp33_ASAP7_75t_R n_10878 (.A1(n_10680_o_0),
    .A2(n_10725_o_0),
    .B(n_10638_o_0),
    .Y(n_10878_o_0));
 INVx1_ASAP7_75t_R n_10879 (.A(n_10718_o_0),
    .Y(n_10879_o_0));
 AOI21xp33_ASAP7_75t_R n_1088 (.A1(n_864_o_0),
    .A2(n_847_o_0),
    .B(n_881_o_0),
    .Y(n_1088_o_0));
 NAND3xp33_ASAP7_75t_R n_10880 (.A(n_10843_o_0),
    .B(n_10723_o_0),
    .C(n_10604_o_0),
    .Y(n_10880_o_0));
 OAI31xp33_ASAP7_75t_R n_10881 (.A1(n_10655_o_0),
    .A2(n_10879_o_0),
    .A3(n_10790_o_0),
    .B(n_10880_o_0),
    .Y(n_10881_o_0));
 AOI21xp33_ASAP7_75t_R n_10882 (.A1(n_10624_o_0),
    .A2(n_10881_o_0),
    .B(n_10648_o_0),
    .Y(n_10882_o_0));
 OAI21xp33_ASAP7_75t_R n_10883 (.A1(n_10611_o_0),
    .A2(n_10878_o_0),
    .B(n_10882_o_0),
    .Y(n_10883_o_0));
 AOI21xp33_ASAP7_75t_R n_10884 (.A1(n_10591_o_0),
    .A2(n_10618_o_0),
    .B(n_10620_o_0),
    .Y(n_10884_o_0));
 OAI21xp33_ASAP7_75t_R n_10885 (.A1(net6),
    .A2(n_10825_o_0),
    .B(n_10884_o_0),
    .Y(n_10885_o_0));
 OAI31xp33_ASAP7_75t_R n_10886 (.A1(n_10655_o_0),
    .A2(n_10677_o_0),
    .A3(n_10663_o_0),
    .B(n_10885_o_0),
    .Y(n_10886_o_0));
 AOI211xp5_ASAP7_75t_R n_10887 (.A1(n_10886_o_0),
    .A2(n_10641_o_0),
    .B(n_10701_o_0),
    .C(n_10832_o_0),
    .Y(n_10887_o_0));
 INVx1_ASAP7_75t_R n_10888 (.A(n_10887_o_0),
    .Y(n_10888_o_0));
 NOR2xp33_ASAP7_75t_R n_10889 (.A(n_10580_o_0),
    .B(n_10643_o_0),
    .Y(n_10889_o_0));
 OAI311xp33_ASAP7_75t_R n_1089 (.A1(n_859_o_0),
    .A2(n_877_o_0),
    .A3(n_1088_o_0),
    .B1(n_983_o_0),
    .C1(n_985_o_0),
    .Y(n_1089_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_10890 (.A1(n_10653_o_0),
    .A2(n_10766_o_0),
    .B(n_10636_o_0),
    .C(n_10621_o_0),
    .D(n_10889_o_0),
    .Y(n_10890_o_0));
 AOI211xp5_ASAP7_75t_R n_10891 (.A1(n_10653_o_0),
    .A2(n_10766_o_0),
    .B(n_10812_o_0),
    .C(n_10632_o_0),
    .Y(n_10891_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10892 (.A1(n_10890_o_0),
    .A2(n_10648_o_0),
    .B(n_10891_o_0),
    .C(n_10700_o_0),
    .Y(n_10892_o_0));
 NAND2xp33_ASAP7_75t_R n_10893 (.A(n_10700_o_0),
    .B(n_10625_o_0),
    .Y(n_10893_o_0));
 INVx1_ASAP7_75t_R n_10894 (.A(n_10595_o_0),
    .Y(n_10894_o_0));
 AOI31xp33_ASAP7_75t_R n_10895 (.A1(net6),
    .A2(n_10825_o_0),
    .A3(n_10655_o_0),
    .B(n_10611_o_0),
    .Y(n_10895_o_0));
 OAI31xp33_ASAP7_75t_R n_10896 (.A1(n_10655_o_0),
    .A2(n_10894_o_0),
    .A3(n_10592_o_0),
    .B(n_10895_o_0),
    .Y(n_10896_o_0));
 NOR2xp33_ASAP7_75t_R n_10897 (.A(n_10701_o_0),
    .B(n_10611_o_0),
    .Y(n_10897_o_0));
 INVx1_ASAP7_75t_R n_10898 (.A(n_10897_o_0),
    .Y(n_10898_o_0));
 OAI211xp5_ASAP7_75t_R n_10899 (.A1(net43),
    .A2(n_10635_o_0),
    .B(n_10718_o_0),
    .C(n_10655_o_0),
    .Y(n_10899_o_0));
 NOR2xp33_ASAP7_75t_R n_1090 (.A(net42),
    .B(n_1089_o_0),
    .Y(n_1090_o_0));
 OAI31xp33_ASAP7_75t_R n_10900 (.A1(n_10655_o_0),
    .A2(n_10664_o_0),
    .A3(n_10790_o_0),
    .B(n_10899_o_0),
    .Y(n_10900_o_0));
 AOI22xp33_ASAP7_75t_R n_10901 (.A1(n_10896_o_0),
    .A2(n_10898_o_0),
    .B1(n_10900_o_0),
    .B2(n_10648_o_0),
    .Y(n_10901_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10902 (.A1(n_10625_o_0),
    .A2(n_10892_o_0),
    .B(n_10893_o_0),
    .C(n_10901_o_0),
    .Y(n_10902_o_0));
 AOI31xp33_ASAP7_75t_R n_10903 (.A1(n_10555_o_0),
    .A2(n_10883_o_0),
    .A3(n_10888_o_0),
    .B(n_10902_o_0),
    .Y(n_10903_o_0));
 INVx1_ASAP7_75t_R n_10904 (.A(n_10767_o_0),
    .Y(n_10904_o_0));
 INVx1_ASAP7_75t_R n_10905 (.A(n_10843_o_0),
    .Y(n_10905_o_0));
 OAI21xp33_ASAP7_75t_R n_10906 (.A1(n_10757_o_0),
    .A2(n_10905_o_0),
    .B(n_10855_o_0),
    .Y(n_10906_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10907 (.A1(net43),
    .A2(n_10614_o_0),
    .B(n_10904_o_0),
    .C(n_10906_o_0),
    .Y(n_10907_o_0));
 NOR2xp33_ASAP7_75t_R n_10908 (.A(n_10567_o_0),
    .B(n_10618_o_0),
    .Y(n_10908_o_0));
 AOI311xp33_ASAP7_75t_R n_10909 (.A1(net12),
    .A2(n_10653_o_0),
    .A3(n_10766_o_0),
    .B(n_10655_o_0),
    .C(n_10908_o_0),
    .Y(n_10909_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1091 (.A1(net16),
    .A2(n_1087_o_0),
    .B(n_1090_o_0),
    .C(n_903_o_0),
    .Y(n_1091_o_0));
 AOI31xp33_ASAP7_75t_R n_10910 (.A1(n_10604_o_0),
    .A2(n_10644_o_0),
    .A3(n_10704_o_0),
    .B(n_10909_o_0),
    .Y(n_10910_o_0));
 OAI21xp33_ASAP7_75t_R n_10911 (.A1(n_10788_o_0),
    .A2(n_10790_o_0),
    .B(n_10623_o_0),
    .Y(n_10911_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10912 (.A1(n_10726_o_0),
    .A2(n_10761_o_0),
    .B(n_10741_o_0),
    .C(n_10624_o_0),
    .Y(n_10912_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10913 (.A1(n_10726_o_0),
    .A2(n_10722_o_0),
    .B(n_10911_o_0),
    .C(n_10912_o_0),
    .Y(n_10913_o_0));
 OAI32xp33_ASAP7_75t_R n_10914 (.A1(n_10611_o_0),
    .A2(n_10910_o_0),
    .A3(n_10632_o_0),
    .B1(n_10913_o_0),
    .B2(n_10701_o_0),
    .Y(n_10914_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10915 (.A1(n_10766_o_0),
    .A2(n_10653_o_0),
    .B(n_10580_o_0),
    .C(n_10639_o_0),
    .Y(n_10915_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10916 (.A1(n_10594_o_0),
    .A2(net43),
    .B(n_10915_o_0),
    .C(n_10724_o_0),
    .Y(n_10916_o_0));
 AOI211xp5_ASAP7_75t_R n_10917 (.A1(net6),
    .A2(n_10825_o_0),
    .B(n_10711_o_0),
    .C(n_10639_o_0),
    .Y(n_10917_o_0));
 NAND3xp33_ASAP7_75t_R n_10918 (.A(n_10766_o_0),
    .B(n_10653_o_0),
    .C(net43),
    .Y(n_10918_o_0));
 AOI21xp33_ASAP7_75t_R n_10919 (.A1(n_10918_o_0),
    .A2(n_10777_o_0),
    .B(n_10655_o_0),
    .Y(n_10919_o_0));
 AOI21xp33_ASAP7_75t_R n_1092 (.A1(n_1084_o_0),
    .A2(n_1091_o_0),
    .B(n_930_o_0),
    .Y(n_1092_o_0));
 OAI211xp5_ASAP7_75t_R n_10920 (.A1(n_10917_o_0),
    .A2(n_10919_o_0),
    .B(n_10641_o_0),
    .C(n_10701_o_0),
    .Y(n_10920_o_0));
 AOI31xp33_ASAP7_75t_R n_10921 (.A1(n_10620_o_0),
    .A2(n_10595_o_0),
    .A3(n_10781_o_0),
    .B(n_10641_o_0),
    .Y(n_10921_o_0));
 INVx1_ASAP7_75t_R n_10922 (.A(n_10921_o_0),
    .Y(n_10922_o_0));
 AOI21xp33_ASAP7_75t_R n_10923 (.A1(n_10722_o_0),
    .A2(n_10726_o_0),
    .B(n_10624_o_0),
    .Y(n_10923_o_0));
 OAI21xp33_ASAP7_75t_R n_10924 (.A1(n_10639_o_0),
    .A2(n_10711_o_0),
    .B(n_10923_o_0),
    .Y(n_10924_o_0));
 OAI211xp5_ASAP7_75t_R n_10925 (.A1(n_10922_o_0),
    .A2(n_10779_o_0),
    .B(n_10648_o_0),
    .C(n_10924_o_0),
    .Y(n_10925_o_0));
 OAI311xp33_ASAP7_75t_R n_10926 (.A1(n_10648_o_0),
    .A2(n_10641_o_0),
    .A3(n_10916_o_0),
    .B1(n_10920_o_0),
    .C1(n_10925_o_0),
    .Y(n_10926_o_0));
 OAI321xp33_ASAP7_75t_R n_10927 (.A1(n_10555_o_0),
    .A2(n_10907_o_0),
    .A3(n_10914_o_0),
    .B1(n_10926_o_0),
    .B2(n_10700_o_0),
    .C(n_10837_o_0),
    .Y(n_10927_o_0));
 OAI21xp33_ASAP7_75t_R n_10928 (.A1(n_10697_o_0),
    .A2(n_10903_o_0),
    .B(n_10927_o_0),
    .Y(n_10928_o_0));
 AOI21xp33_ASAP7_75t_R n_10929 (.A1(n_10852_o_0),
    .A2(n_10722_o_0),
    .B(n_10604_o_0),
    .Y(n_10929_o_0));
 INVx1_ASAP7_75t_R n_1093 (.A(n_989_o_0),
    .Y(n_1093_o_0));
 AOI21xp33_ASAP7_75t_R n_10930 (.A1(n_10595_o_0),
    .A2(n_10792_o_0),
    .B(n_10620_o_0),
    .Y(n_10930_o_0));
 AO21x1_ASAP7_75t_R n_10931 (.A1(n_10724_o_0),
    .A2(n_10686_o_0),
    .B(n_10611_o_0),
    .Y(n_10931_o_0));
 OAI31xp33_ASAP7_75t_R n_10932 (.A1(n_10623_o_0),
    .A2(n_10929_o_0),
    .A3(n_10930_o_0),
    .B(n_10931_o_0),
    .Y(n_10932_o_0));
 AND3x1_ASAP7_75t_R n_10933 (.A(n_10595_o_0),
    .B(n_10764_o_0),
    .C(n_10604_o_0),
    .Y(n_10933_o_0));
 AOI31xp33_ASAP7_75t_R n_10934 (.A1(net12),
    .A2(n_10620_o_0),
    .A3(n_10722_o_0),
    .B(n_10933_o_0),
    .Y(n_10934_o_0));
 AOI31xp33_ASAP7_75t_R n_10935 (.A1(n_10591_o_0),
    .A2(n_10639_o_0),
    .A3(n_10567_o_0),
    .B(n_10611_o_0),
    .Y(n_10935_o_0));
 NOR3xp33_ASAP7_75t_R n_10936 (.A(n_10654_o_0),
    .B(n_10620_o_0),
    .C(net6),
    .Y(n_10936_o_0));
 INVx1_ASAP7_75t_R n_10937 (.A(n_10936_o_0),
    .Y(n_10937_o_0));
 AOI21xp33_ASAP7_75t_R n_10938 (.A1(n_10935_o_0),
    .A2(n_10937_o_0),
    .B(n_10648_o_0),
    .Y(n_10938_o_0));
 OAI21xp33_ASAP7_75t_R n_10939 (.A1(n_10623_o_0),
    .A2(n_10934_o_0),
    .B(n_10938_o_0),
    .Y(n_10939_o_0));
 NAND3xp33_ASAP7_75t_R n_1094 (.A(n_1093_o_0),
    .B(n_909_o_0),
    .C(n_878_o_0),
    .Y(n_1094_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10940 (.A1(n_10633_o_0),
    .A2(n_10932_o_0),
    .B(n_10939_o_0),
    .C(n_10837_o_0),
    .Y(n_10940_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10941 (.A1(net12),
    .A2(n_10815_o_0),
    .B(n_10817_o_0),
    .C(n_10624_o_0),
    .Y(n_10941_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10942 (.A1(net12),
    .A2(n_10661_o_0),
    .B(n_10669_o_0),
    .C(n_10604_o_0),
    .Y(n_10942_o_0));
 OAI21xp33_ASAP7_75t_R n_10943 (.A1(n_10620_o_0),
    .A2(n_10669_o_0),
    .B(n_10624_o_0),
    .Y(n_10943_o_0));
 OAI31xp33_ASAP7_75t_R n_10944 (.A1(n_10936_o_0),
    .A2(n_10942_o_0),
    .A3(n_10943_o_0),
    .B(n_10633_o_0),
    .Y(n_10944_o_0));
 OAI211xp5_ASAP7_75t_R n_10945 (.A1(n_10683_o_0),
    .A2(net43),
    .B(n_10718_o_0),
    .C(n_10639_o_0),
    .Y(n_10945_o_0));
 OAI31xp33_ASAP7_75t_R n_10946 (.A1(n_10639_o_0),
    .A2(n_10838_o_0),
    .A3(n_10908_o_0),
    .B(n_10945_o_0),
    .Y(n_10946_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10947 (.A1(net12),
    .A2(n_10591_o_0),
    .B(n_10567_o_0),
    .C(n_10604_o_0),
    .Y(n_10947_o_0));
 AOI31xp33_ASAP7_75t_R n_10948 (.A1(n_10947_o_0),
    .A2(n_10645_o_0),
    .A3(n_10623_o_0),
    .B(n_10701_o_0),
    .Y(n_10948_o_0));
 OAI21xp33_ASAP7_75t_R n_10949 (.A1(n_10641_o_0),
    .A2(n_10946_o_0),
    .B(n_10948_o_0),
    .Y(n_10949_o_0));
 AOI21xp33_ASAP7_75t_R n_1095 (.A1(n_877_o_0),
    .A2(n_956_o_0),
    .B(n_904_o_0),
    .Y(n_1095_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10950 (.A1(n_10941_o_0),
    .A2(n_10605_o_0),
    .B(n_10944_o_0),
    .C(n_10949_o_0),
    .Y(n_10950_o_0));
 NOR2xp33_ASAP7_75t_R n_10951 (.A(n_10696_o_0),
    .B(n_10950_o_0),
    .Y(n_10951_o_0));
 AOI21xp33_ASAP7_75t_R n_10952 (.A1(n_10620_o_0),
    .A2(n_10818_o_0),
    .B(n_10782_o_0),
    .Y(n_10952_o_0));
 AOI211xp5_ASAP7_75t_R n_10953 (.A1(n_10918_o_0),
    .A2(n_10857_o_0),
    .B(n_10665_o_0),
    .C(n_10611_o_0),
    .Y(n_10953_o_0));
 AOI211xp5_ASAP7_75t_R n_10954 (.A1(n_10611_o_0),
    .A2(n_10952_o_0),
    .B(n_10953_o_0),
    .C(n_10632_o_0),
    .Y(n_10954_o_0));
 AOI21xp33_ASAP7_75t_R n_10955 (.A1(n_10718_o_0),
    .A2(n_10726_o_0),
    .B(n_10670_o_0),
    .Y(n_10955_o_0));
 NAND3xp33_ASAP7_75t_R n_10956 (.A(n_10620_o_0),
    .B(n_10643_o_0),
    .C(net43),
    .Y(n_10956_o_0));
 OAI211xp5_ASAP7_75t_R n_10957 (.A1(n_10740_o_0),
    .A2(n_10655_o_0),
    .B(n_10956_o_0),
    .C(n_10801_o_0),
    .Y(n_10957_o_0));
 OAI21xp33_ASAP7_75t_R n_10958 (.A1(n_10641_o_0),
    .A2(n_10957_o_0),
    .B(n_10648_o_0),
    .Y(n_10958_o_0));
 AOI21xp33_ASAP7_75t_R n_10959 (.A1(n_10623_o_0),
    .A2(n_10955_o_0),
    .B(n_10958_o_0),
    .Y(n_10959_o_0));
 OAI21xp33_ASAP7_75t_R n_1096 (.A1(n_935_o_0),
    .A2(net32),
    .B(n_893_o_0),
    .Y(n_1096_o_0));
 OAI21xp33_ASAP7_75t_R n_10960 (.A1(n_10635_o_0),
    .A2(net6),
    .B(n_10643_o_0),
    .Y(n_10960_o_0));
 AOI211xp5_ASAP7_75t_R n_10961 (.A1(n_10960_o_0),
    .A2(n_10604_o_0),
    .B(n_10929_o_0),
    .C(n_10641_o_0),
    .Y(n_10961_o_0));
 INVx1_ASAP7_75t_R n_10962 (.A(n_10847_o_0),
    .Y(n_10962_o_0));
 AOI211xp5_ASAP7_75t_R n_10963 (.A1(n_10726_o_0),
    .A2(n_10761_o_0),
    .B(n_10962_o_0),
    .C(n_10624_o_0),
    .Y(n_10963_o_0));
 OAI21xp33_ASAP7_75t_R n_10964 (.A1(n_10639_o_0),
    .A2(n_10894_o_0),
    .B(n_10611_o_0),
    .Y(n_10964_o_0));
 OAI21xp33_ASAP7_75t_R n_10965 (.A1(n_10618_o_0),
    .A2(n_10643_o_0),
    .B(n_10604_o_0),
    .Y(n_10965_o_0));
 AOI21xp33_ASAP7_75t_R n_10966 (.A1(n_10731_o_0),
    .A2(n_10803_o_0),
    .B(n_10624_o_0),
    .Y(n_10966_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10967 (.A1(n_10965_o_0),
    .A2(n_10592_o_0),
    .B(n_10966_o_0),
    .C(n_10632_o_0),
    .Y(n_10967_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10968 (.A1(net12),
    .A2(n_10614_o_0),
    .B(n_10964_o_0),
    .C(n_10967_o_0),
    .Y(n_10968_o_0));
 OAI31xp33_ASAP7_75t_R n_10969 (.A1(n_10701_o_0),
    .A2(n_10961_o_0),
    .A3(n_10963_o_0),
    .B(n_10968_o_0),
    .Y(n_10969_o_0));
 OAI21xp33_ASAP7_75t_R n_1097 (.A1(n_878_o_0),
    .A2(n_1093_o_0),
    .B(n_1096_o_0),
    .Y(n_1097_o_0));
 OAI321xp33_ASAP7_75t_R n_10970 (.A1(n_10837_o_0),
    .A2(n_10954_o_0),
    .A3(n_10959_o_0),
    .B1(n_10969_o_0),
    .B2(n_10696_o_0),
    .C(n_10555_o_0),
    .Y(n_10970_o_0));
 OAI31xp33_ASAP7_75t_R n_10971 (.A1(n_10796_o_0),
    .A2(n_10940_o_0),
    .A3(n_10951_o_0),
    .B(n_10970_o_0),
    .Y(n_10971_o_0));
 AOI21xp33_ASAP7_75t_R n_10972 (.A1(n_10567_o_0),
    .A2(n_10655_o_0),
    .B(n_10929_o_0),
    .Y(n_10972_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10973 (.A1(n_10663_o_0),
    .A2(n_10677_o_0),
    .B(n_10604_o_0),
    .C(n_10641_o_0),
    .Y(n_10973_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10974 (.A1(n_10591_o_0),
    .A2(n_10567_o_0),
    .B(n_10713_o_0),
    .C(n_10973_o_0),
    .Y(n_10974_o_0));
 OAI211xp5_ASAP7_75t_R n_10975 (.A1(n_10624_o_0),
    .A2(n_10972_o_0),
    .B(n_10974_o_0),
    .C(n_10633_o_0),
    .Y(n_10975_o_0));
 OAI211xp5_ASAP7_75t_R n_10976 (.A1(net12),
    .A2(n_10635_o_0),
    .B(n_10643_o_0),
    .C(n_10639_o_0),
    .Y(n_10976_o_0));
 NOR2xp33_ASAP7_75t_R n_10977 (.A(n_10701_o_0),
    .B(n_10623_o_0),
    .Y(n_10977_o_0));
 NAND3xp33_ASAP7_75t_R n_10978 (.A(n_10567_o_0),
    .B(net43),
    .C(n_10591_o_0),
    .Y(n_10978_o_0));
 AOI22xp33_ASAP7_75t_R n_10979 (.A1(n_10717_o_0),
    .A2(n_10818_o_0),
    .B1(n_10620_o_0),
    .B2(n_10978_o_0),
    .Y(n_10979_o_0));
 OAI21xp33_ASAP7_75t_R n_1098 (.A1(n_903_o_0),
    .A2(n_1097_o_0),
    .B(net15),
    .Y(n_1098_o_0));
 NOR2xp33_ASAP7_75t_R n_10980 (.A(n_10898_o_0),
    .B(n_10979_o_0),
    .Y(n_10980_o_0));
 AOI31xp33_ASAP7_75t_R n_10981 (.A1(n_10937_o_0),
    .A2(n_10976_o_0),
    .A3(n_10977_o_0),
    .B(n_10980_o_0),
    .Y(n_10981_o_0));
 AOI21xp33_ASAP7_75t_R n_10982 (.A1(n_10975_o_0),
    .A2(n_10981_o_0),
    .B(n_10796_o_0),
    .Y(n_10982_o_0));
 NAND3xp33_ASAP7_75t_R n_10983 (.A(n_10772_o_0),
    .B(n_10718_o_0),
    .C(n_10604_o_0),
    .Y(n_10983_o_0));
 AOI211xp5_ASAP7_75t_R n_10984 (.A1(n_10643_o_0),
    .A2(net43),
    .B(n_10639_o_0),
    .C(n_10591_o_0),
    .Y(n_10984_o_0));
 AOI311xp33_ASAP7_75t_R n_10985 (.A1(n_10620_o_0),
    .A2(n_10593_o_0),
    .A3(n_10595_o_0),
    .B(n_10641_o_0),
    .C(n_10984_o_0),
    .Y(n_10985_o_0));
 AOI31xp33_ASAP7_75t_R n_10986 (.A1(n_10956_o_0),
    .A2(n_10983_o_0),
    .A3(n_10617_o_0),
    .B(n_10985_o_0),
    .Y(n_10986_o_0));
 INVx1_ASAP7_75t_R n_10987 (.A(n_10915_o_0),
    .Y(n_10987_o_0));
 AOI21xp33_ASAP7_75t_R n_10988 (.A1(n_10702_o_0),
    .A2(n_10669_o_0),
    .B(n_10620_o_0),
    .Y(n_10988_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_10989 (.A1(n_10643_o_0),
    .A2(n_10591_o_0),
    .B(net43),
    .C(n_10623_o_0),
    .Y(n_10989_o_0));
 AOI21xp33_ASAP7_75t_R n_1099 (.A1(n_1094_o_0),
    .A2(n_1095_o_0),
    .B(n_1098_o_0),
    .Y(n_1099_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_10990 (.A1(n_10661_o_0),
    .A2(net12),
    .B(n_10604_o_0),
    .C(n_10989_o_0),
    .Y(n_10990_o_0));
 OAI31xp33_ASAP7_75t_R n_10991 (.A1(n_10611_o_0),
    .A2(n_10987_o_0),
    .A3(n_10988_o_0),
    .B(n_10990_o_0),
    .Y(n_10991_o_0));
 OAI21xp33_ASAP7_75t_R n_10992 (.A1(n_10633_o_0),
    .A2(n_10991_o_0),
    .B(n_10555_o_0),
    .Y(n_10992_o_0));
 AOI21xp33_ASAP7_75t_R n_10993 (.A1(n_10633_o_0),
    .A2(n_10986_o_0),
    .B(n_10992_o_0),
    .Y(n_10993_o_0));
 NOR2xp33_ASAP7_75t_R n_10994 (.A(n_10805_o_0),
    .B(n_10806_o_0),
    .Y(n_10994_o_0));
 INVx1_ASAP7_75t_R n_10995 (.A(n_10884_o_0),
    .Y(n_10995_o_0));
 OAI211xp5_ASAP7_75t_R n_10996 (.A1(n_10994_o_0),
    .A2(n_10655_o_0),
    .B(n_10995_o_0),
    .C(n_10701_o_0),
    .Y(n_10996_o_0));
 AOI21xp33_ASAP7_75t_R n_10997 (.A1(n_10604_o_0),
    .A2(n_10594_o_0),
    .B(n_10633_o_0),
    .Y(n_10997_o_0));
 OAI21xp33_ASAP7_75t_R n_10998 (.A1(n_10655_o_0),
    .A2(n_10663_o_0),
    .B(n_10997_o_0),
    .Y(n_10998_o_0));
 AND3x1_ASAP7_75t_R n_10999 (.A(n_10996_o_0),
    .B(n_10998_o_0),
    .C(n_10641_o_0),
    .Y(n_10999_o_0));
 OAI311xp33_ASAP7_75t_R n_1100 (.A1(net32),
    .A2(n_1028_o_0),
    .A3(n_917_o_0),
    .B1(n_990_o_0),
    .C1(n_878_o_0),
    .Y(n_1100_o_0));
 INVx1_ASAP7_75t_R n_11000 (.A(n_10977_o_0),
    .Y(n_11000_o_0));
 AOI211xp5_ASAP7_75t_R n_11001 (.A1(net6),
    .A2(n_10654_o_0),
    .B(n_10677_o_0),
    .C(n_10639_o_0),
    .Y(n_11001_o_0));
 AOI31xp33_ASAP7_75t_R n_11002 (.A1(n_10620_o_0),
    .A2(n_10718_o_0),
    .A3(n_10781_o_0),
    .B(n_11001_o_0),
    .Y(n_11002_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11003 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(net43),
    .C(n_10620_o_0),
    .Y(n_11003_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11004 (.A1(n_11003_o_0),
    .A2(n_10662_o_0),
    .B(n_10855_o_0),
    .C(n_10796_o_0),
    .Y(n_11004_o_0));
 OAI21xp33_ASAP7_75t_R n_11005 (.A1(n_11000_o_0),
    .A2(n_11002_o_0),
    .B(n_11004_o_0),
    .Y(n_11005_o_0));
 AND3x1_ASAP7_75t_R n_11006 (.A(n_10595_o_0),
    .B(n_10764_o_0),
    .C(n_10620_o_0),
    .Y(n_11006_o_0));
 AOI21xp33_ASAP7_75t_R n_11007 (.A1(n_10717_o_0),
    .A2(n_10710_o_0),
    .B(n_11006_o_0),
    .Y(n_11007_o_0));
 OAI31xp33_ASAP7_75t_R n_11008 (.A1(n_10655_o_0),
    .A2(n_10879_o_0),
    .A3(n_10663_o_0),
    .B(n_10632_o_0),
    .Y(n_11008_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11009 (.A1(n_10594_o_0),
    .A2(n_10670_o_0),
    .B(n_11008_o_0),
    .C(n_10624_o_0),
    .Y(n_11009_o_0));
 OAI31xp33_ASAP7_75t_R n_1101 (.A1(n_878_o_0),
    .A2(n_915_o_0),
    .A3(n_989_o_0),
    .B(n_1100_o_0),
    .Y(n_1101_o_0));
 NAND2xp33_ASAP7_75t_R n_11010 (.A(n_10644_o_0),
    .B(n_10803_o_0),
    .Y(n_11010_o_0));
 OAI31xp33_ASAP7_75t_R n_11011 (.A1(n_10639_o_0),
    .A2(n_10664_o_0),
    .A3(n_10663_o_0),
    .B(n_11010_o_0),
    .Y(n_11011_o_0));
 NAND2xp33_ASAP7_75t_R n_11012 (.A(n_10591_o_0),
    .B(n_10604_o_0),
    .Y(n_11012_o_0));
 AOI211xp5_ASAP7_75t_R n_11013 (.A1(n_10727_o_0),
    .A2(n_11012_o_0),
    .B(n_10611_o_0),
    .C(n_10632_o_0),
    .Y(n_11013_o_0));
 AOI21xp33_ASAP7_75t_R n_11014 (.A1(n_10897_o_0),
    .A2(n_11011_o_0),
    .B(n_11013_o_0),
    .Y(n_11014_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11015 (.A1(n_10701_o_0),
    .A2(n_11007_o_0),
    .B(n_11009_o_0),
    .C(n_11014_o_0),
    .Y(n_11015_o_0));
 OAI221xp5_ASAP7_75t_R n_11016 (.A1(n_10999_o_0),
    .A2(n_11005_o_0),
    .B1(n_10700_o_0),
    .B2(n_11015_o_0),
    .C(n_10696_o_0),
    .Y(n_11016_o_0));
 OAI31xp33_ASAP7_75t_R n_11017 (.A1(n_10754_o_0),
    .A2(n_10982_o_0),
    .A3(n_10993_o_0),
    .B(n_11016_o_0),
    .Y(n_11017_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11018 (.A1(n_10639_o_0),
    .A2(n_10649_o_0),
    .B(n_10703_o_0),
    .C(n_10632_o_0),
    .Y(n_11018_o_0));
 OAI21xp33_ASAP7_75t_R n_11019 (.A1(n_10604_o_0),
    .A2(n_10746_o_0),
    .B(n_11018_o_0),
    .Y(n_11019_o_0));
 OAI21xp33_ASAP7_75t_R n_1102 (.A1(n_907_o_0),
    .A2(n_887_o_0),
    .B(n_878_o_0),
    .Y(n_1102_o_0));
 OAI21xp33_ASAP7_75t_R n_11020 (.A1(n_10635_o_0),
    .A2(n_10580_o_0),
    .B(n_10567_o_0),
    .Y(n_11020_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11021 (.A1(n_11020_o_0),
    .A2(n_10604_o_0),
    .B(n_10742_o_0),
    .C(n_10648_o_0),
    .Y(n_11021_o_0));
 NAND3xp33_ASAP7_75t_R n_11022 (.A(n_11019_o_0),
    .B(n_11021_o_0),
    .C(n_10611_o_0),
    .Y(n_11022_o_0));
 AOI211xp5_ASAP7_75t_R n_11023 (.A1(n_10815_o_0),
    .A2(net6),
    .B(n_10655_o_0),
    .C(n_10685_o_0),
    .Y(n_11023_o_0));
 AOI31xp33_ASAP7_75t_R n_11024 (.A1(n_10604_o_0),
    .A2(n_10764_o_0),
    .A3(n_10710_o_0),
    .B(n_11023_o_0),
    .Y(n_11024_o_0));
 INVx1_ASAP7_75t_R n_11025 (.A(n_10679_o_0),
    .Y(n_11025_o_0));
 OAI211xp5_ASAP7_75t_R n_11026 (.A1(n_10676_o_0),
    .A2(n_10643_o_0),
    .B(n_10604_o_0),
    .C(n_10723_o_0),
    .Y(n_11026_o_0));
 OAI31xp33_ASAP7_75t_R n_11027 (.A1(n_10655_o_0),
    .A2(n_11025_o_0),
    .A3(n_10870_o_0),
    .B(n_11026_o_0),
    .Y(n_11027_o_0));
 AOI21xp33_ASAP7_75t_R n_11028 (.A1(n_10648_o_0),
    .A2(n_11027_o_0),
    .B(n_10624_o_0),
    .Y(n_11028_o_0));
 OAI21xp33_ASAP7_75t_R n_11029 (.A1(n_10632_o_0),
    .A2(n_11024_o_0),
    .B(n_11028_o_0),
    .Y(n_11029_o_0));
 OAI21xp33_ASAP7_75t_R n_1103 (.A1(n_989_o_0),
    .A2(n_991_o_0),
    .B(n_1102_o_0),
    .Y(n_1103_o_0));
 AOI211xp5_ASAP7_75t_R n_11030 (.A1(n_10635_o_0),
    .A2(n_10567_o_0),
    .B(n_10908_o_0),
    .C(n_10639_o_0),
    .Y(n_11030_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11031 (.A1(n_10643_o_0),
    .A2(n_10639_o_0),
    .B(n_11030_o_0),
    .C(n_10701_o_0),
    .Y(n_11031_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11032 (.A1(net12),
    .A2(n_10615_o_0),
    .B(n_10816_o_0),
    .C(n_10632_o_0),
    .Y(n_11032_o_0));
 AOI21xp33_ASAP7_75t_R n_11033 (.A1(n_10595_o_0),
    .A2(n_10817_o_0),
    .B(n_11032_o_0),
    .Y(n_11033_o_0));
 OAI21xp33_ASAP7_75t_R n_11034 (.A1(net6),
    .A2(n_10654_o_0),
    .B(n_10726_o_0),
    .Y(n_11034_o_0));
 OAI31xp33_ASAP7_75t_R n_11035 (.A1(n_10591_o_0),
    .A2(n_10639_o_0),
    .A3(net6),
    .B(n_11034_o_0),
    .Y(n_11035_o_0));
 AOI22xp33_ASAP7_75t_R n_11036 (.A1(n_10670_o_0),
    .A2(n_10614_o_0),
    .B1(n_10620_o_0),
    .B2(n_10739_o_0),
    .Y(n_11036_o_0));
 OAI221xp5_ASAP7_75t_R n_11037 (.A1(n_10620_o_0),
    .A2(n_10669_o_0),
    .B1(n_10632_o_0),
    .B2(n_11036_o_0),
    .C(n_10624_o_0),
    .Y(n_11037_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11038 (.A1(n_10632_o_0),
    .A2(n_11035_o_0),
    .B(n_11037_o_0),
    .C(n_10796_o_0),
    .Y(n_11038_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11039 (.A1(n_10701_o_0),
    .A2(n_11031_o_0),
    .B(n_11033_o_0),
    .C(n_10623_o_0),
    .D(n_11038_o_0),
    .Y(n_11039_o_0));
 OAI21xp33_ASAP7_75t_R n_1104 (.A1(n_903_o_0),
    .A2(n_1103_o_0),
    .B(net16),
    .Y(n_1104_o_0));
 AOI31xp33_ASAP7_75t_R n_11040 (.A1(n_10700_o_0),
    .A2(n_11022_o_0),
    .A3(n_11029_o_0),
    .B(n_11039_o_0),
    .Y(n_11040_o_0));
 XOR2xp5_ASAP7_75t_R n_11041 (.A(net43),
    .B(n_10643_o_0),
    .Y(n_11041_o_0));
 AOI211xp5_ASAP7_75t_R n_11042 (.A1(n_10604_o_0),
    .A2(n_11041_o_0),
    .B(n_11006_o_0),
    .C(n_10624_o_0),
    .Y(n_11042_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11043 (.A1(n_10717_o_0),
    .A2(n_10978_o_0),
    .B(n_10811_o_0),
    .C(n_10855_o_0),
    .Y(n_11043_o_0));
 OAI321xp33_ASAP7_75t_R n_11044 (.A1(n_11000_o_0),
    .A2(n_10933_o_0),
    .A3(n_10622_o_0),
    .B1(n_10860_o_0),
    .B2(n_10898_o_0),
    .C(n_11043_o_0),
    .Y(n_11044_o_0));
 AOI21xp33_ASAP7_75t_R n_11045 (.A1(n_10701_o_0),
    .A2(n_11042_o_0),
    .B(n_11044_o_0),
    .Y(n_11045_o_0));
 AOI32xp33_ASAP7_75t_R n_11046 (.A1(n_10604_o_0),
    .A2(n_10702_o_0),
    .A3(n_10669_o_0),
    .B1(n_10781_o_0),
    .B2(n_10620_o_0),
    .Y(n_11046_o_0));
 AOI21xp33_ASAP7_75t_R n_11047 (.A1(n_10762_o_0),
    .A2(n_10715_o_0),
    .B(n_10701_o_0),
    .Y(n_11047_o_0));
 OAI21xp33_ASAP7_75t_R n_11048 (.A1(n_10624_o_0),
    .A2(n_11046_o_0),
    .B(n_11047_o_0),
    .Y(n_11048_o_0));
 OAI21xp33_ASAP7_75t_R n_11049 (.A1(n_10635_o_0),
    .A2(net6),
    .B(n_10623_o_0),
    .Y(n_11049_o_0));
 AOI21xp33_ASAP7_75t_R n_1105 (.A1(n_903_o_0),
    .A2(n_1101_o_0),
    .B(n_1104_o_0),
    .Y(n_1105_o_0));
 AOI21xp33_ASAP7_75t_R n_11050 (.A1(n_10604_o_0),
    .A2(n_10725_o_0),
    .B(n_10817_o_0),
    .Y(n_11050_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11051 (.A1(n_10591_o_0),
    .A2(net43),
    .B(n_11050_o_0),
    .C(n_10611_o_0),
    .D(n_10632_o_0),
    .Y(n_11051_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11052 (.A1(n_10643_o_0),
    .A2(n_11012_o_0),
    .B(n_11049_o_0),
    .C(n_11051_o_0),
    .Y(n_11052_o_0));
 AOI31xp33_ASAP7_75t_R n_11053 (.A1(n_10796_o_0),
    .A2(n_11048_o_0),
    .A3(n_11052_o_0),
    .B(n_10697_o_0),
    .Y(n_11053_o_0));
 OAI21xp33_ASAP7_75t_R n_11054 (.A1(n_10555_o_0),
    .A2(n_11045_o_0),
    .B(n_11053_o_0),
    .Y(n_11054_o_0));
 OAI21xp33_ASAP7_75t_R n_11055 (.A1(n_10754_o_0),
    .A2(n_11040_o_0),
    .B(n_11054_o_0),
    .Y(n_11055_o_0));
 AOI21xp33_ASAP7_75t_R n_11056 (.A1(n_10781_o_0),
    .A2(n_10904_o_0),
    .B(n_11000_o_0),
    .Y(n_11056_o_0));
 AOI21xp33_ASAP7_75t_R n_11057 (.A1(n_10591_o_0),
    .A2(n_10567_o_0),
    .B(n_10639_o_0),
    .Y(n_11057_o_0));
 INVx1_ASAP7_75t_R n_11058 (.A(n_11020_o_0),
    .Y(n_11058_o_0));
 OAI211xp5_ASAP7_75t_R n_11059 (.A1(n_10655_o_0),
    .A2(n_11058_o_0),
    .B(n_10801_o_0),
    .C(n_10855_o_0),
    .Y(n_11059_o_0));
 OAI21xp33_ASAP7_75t_R n_1106 (.A1(n_877_o_0),
    .A2(n_989_o_0),
    .B(n_936_o_0),
    .Y(n_1106_o_0));
 NAND3xp33_ASAP7_75t_R n_11060 (.A(n_10655_o_0),
    .B(n_10643_o_0),
    .C(n_10580_o_0),
    .Y(n_11060_o_0));
 OAI311xp33_ASAP7_75t_R n_11061 (.A1(n_10655_o_0),
    .A2(n_10905_o_0),
    .A3(n_11025_o_0),
    .B1(n_11060_o_0),
    .C1(n_10897_o_0),
    .Y(n_11061_o_0));
 OAI311xp33_ASAP7_75t_R n_11062 (.A1(n_10648_o_0),
    .A2(n_10642_o_0),
    .A3(n_11057_o_0),
    .B1(n_11059_o_0),
    .C1(n_11061_o_0),
    .Y(n_11062_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11063 (.A1(net12),
    .A2(n_10643_o_0),
    .B(n_10713_o_0),
    .C(n_11056_o_0),
    .D(n_11062_o_0),
    .Y(n_11063_o_0));
 AOI211xp5_ASAP7_75t_R n_11064 (.A1(n_10639_o_0),
    .A2(n_10683_o_0),
    .B(n_11030_o_0),
    .C(n_10641_o_0),
    .Y(n_11064_o_0));
 AOI211xp5_ASAP7_75t_R n_11065 (.A1(n_10670_o_0),
    .A2(n_10643_o_0),
    .B(n_10642_o_0),
    .C(n_10739_o_0),
    .Y(n_11065_o_0));
 AO21x1_ASAP7_75t_R n_11066 (.A1(n_10729_o_0),
    .A2(net43),
    .B(n_10739_o_0),
    .Y(n_11066_o_0));
 NAND2xp33_ASAP7_75t_R n_11067 (.A(n_10623_o_0),
    .B(n_10655_o_0),
    .Y(n_11067_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11068 (.A1(net43),
    .A2(n_10729_o_0),
    .B(n_10739_o_0),
    .C(n_11067_o_0),
    .Y(n_11068_o_0));
 OAI21xp33_ASAP7_75t_R n_11069 (.A1(n_10623_o_0),
    .A2(n_11066_o_0),
    .B(n_11068_o_0),
    .Y(n_11069_o_0));
 INVx1_ASAP7_75t_R n_1107 (.A(n_861_o_0),
    .Y(n_1107_o_0));
 INVx1_ASAP7_75t_R n_11070 (.A(n_10680_o_0),
    .Y(n_11070_o_0));
 AOI21xp33_ASAP7_75t_R n_11071 (.A1(n_10595_o_0),
    .A2(n_10884_o_0),
    .B(n_10641_o_0),
    .Y(n_11071_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11072 (.A1(n_10591_o_0),
    .A2(n_10567_o_0),
    .B(n_11070_o_0),
    .C(n_11071_o_0),
    .D(n_10632_o_0),
    .Y(n_11072_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11073 (.A1(n_10678_o_0),
    .A2(n_10781_o_0),
    .B(n_11069_o_0),
    .C(n_11072_o_0),
    .Y(n_11073_o_0));
 OAI31xp33_ASAP7_75t_R n_11074 (.A1(n_10701_o_0),
    .A2(n_11064_o_0),
    .A3(n_11065_o_0),
    .B(n_11073_o_0),
    .Y(n_11074_o_0));
 AOI22xp33_ASAP7_75t_R n_11075 (.A1(n_11063_o_0),
    .A2(n_10700_o_0),
    .B1(n_10555_o_0),
    .B2(n_11074_o_0),
    .Y(n_11075_o_0));
 AOI31xp33_ASAP7_75t_R n_11076 (.A1(n_10591_o_0),
    .A2(net43),
    .A3(n_10567_o_0),
    .B(n_10655_o_0),
    .Y(n_11076_o_0));
 AOI22xp33_ASAP7_75t_R n_11077 (.A1(n_10593_o_0),
    .A2(n_10604_o_0),
    .B1(n_11076_o_0),
    .B2(n_10781_o_0),
    .Y(n_11077_o_0));
 OAI211xp5_ASAP7_75t_R n_11078 (.A1(n_10620_o_0),
    .A2(n_10778_o_0),
    .B(n_10915_o_0),
    .C(n_10641_o_0),
    .Y(n_11078_o_0));
 OAI21xp33_ASAP7_75t_R n_11079 (.A1(n_10623_o_0),
    .A2(n_11077_o_0),
    .B(n_11078_o_0),
    .Y(n_11079_o_0));
 AOI21xp33_ASAP7_75t_R n_1108 (.A1(n_1029_o_0),
    .A2(n_937_o_0),
    .B(n_903_o_0),
    .Y(n_1108_o_0));
 AOI21xp33_ASAP7_75t_R n_11080 (.A1(n_10635_o_0),
    .A2(n_10643_o_0),
    .B(n_10889_o_0),
    .Y(n_11080_o_0));
 AOI22xp33_ASAP7_75t_R n_11081 (.A1(n_11080_o_0),
    .A2(n_10604_o_0),
    .B1(n_10764_o_0),
    .B2(n_11076_o_0),
    .Y(n_11081_o_0));
 AOI21xp33_ASAP7_75t_R n_11082 (.A1(n_10635_o_0),
    .A2(n_10620_o_0),
    .B(n_10641_o_0),
    .Y(n_11082_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11083 (.A1(n_10592_o_0),
    .A2(n_10965_o_0),
    .B(n_11082_o_0),
    .C(n_10632_o_0),
    .Y(n_11083_o_0));
 OAI21xp33_ASAP7_75t_R n_11084 (.A1(n_10611_o_0),
    .A2(n_11081_o_0),
    .B(n_11083_o_0),
    .Y(n_11084_o_0));
 OA21x2_ASAP7_75t_R n_11085 (.A1(n_10633_o_0),
    .A2(n_11079_o_0),
    .B(n_11084_o_0),
    .Y(n_11085_o_0));
 NAND2xp33_ASAP7_75t_R n_11086 (.A(n_10639_o_0),
    .B(n_10611_o_0),
    .Y(n_11086_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11087 (.A1(net43),
    .A2(n_10729_o_0),
    .B(n_10739_o_0),
    .C(n_11086_o_0),
    .Y(n_11087_o_0));
 OAI21xp33_ASAP7_75t_R n_11088 (.A1(n_10611_o_0),
    .A2(n_11066_o_0),
    .B(n_11087_o_0),
    .Y(n_11088_o_0));
 AOI31xp33_ASAP7_75t_R n_11089 (.A1(n_10604_o_0),
    .A2(n_10595_o_0),
    .A3(n_10764_o_0),
    .B(n_10817_o_0),
    .Y(n_11089_o_0));
 OAI21xp33_ASAP7_75t_R n_1109 (.A1(n_1107_o_0),
    .A2(n_878_o_0),
    .B(n_1108_o_0),
    .Y(n_1109_o_0));
 NAND2xp33_ASAP7_75t_R n_11090 (.A(n_10623_o_0),
    .B(n_11089_o_0),
    .Y(n_11090_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11091 (.A1(n_10593_o_0),
    .A2(n_10712_o_0),
    .B(n_11088_o_0),
    .C(n_11090_o_0),
    .Y(n_11091_o_0));
 NAND2xp33_ASAP7_75t_R n_11092 (.A(n_10817_o_0),
    .B(n_10595_o_0),
    .Y(n_11092_o_0));
 OAI31xp33_ASAP7_75t_R n_11093 (.A1(n_10639_o_0),
    .A2(n_10592_o_0),
    .A3(n_10908_o_0),
    .B(n_11092_o_0),
    .Y(n_11093_o_0));
 OAI22xp33_ASAP7_75t_R n_11094 (.A1(n_10713_o_0),
    .A2(n_10790_o_0),
    .B1(n_10767_o_0),
    .B2(n_10768_o_0),
    .Y(n_11094_o_0));
 AOI22xp33_ASAP7_75t_R n_11095 (.A1(n_11093_o_0),
    .A2(n_10897_o_0),
    .B1(n_11094_o_0),
    .B2(n_10977_o_0),
    .Y(n_11095_o_0));
 OAI211xp5_ASAP7_75t_R n_11096 (.A1(n_11091_o_0),
    .A2(n_10632_o_0),
    .B(n_10796_o_0),
    .C(n_11095_o_0),
    .Y(n_11096_o_0));
 OAI211xp5_ASAP7_75t_R n_11097 (.A1(n_10555_o_0),
    .A2(n_11085_o_0),
    .B(n_11096_o_0),
    .C(n_10696_o_0),
    .Y(n_11097_o_0));
 OAI21xp33_ASAP7_75t_R n_11098 (.A1(n_10754_o_0),
    .A2(n_11075_o_0),
    .B(n_11097_o_0),
    .Y(n_11098_o_0));
 XOR2xp5_ASAP7_75t_R n_11099 (.A(_01017_),
    .B(_01104_),
    .Y(n_11099_o_0));
 OAI211xp5_ASAP7_75t_R n_1110 (.A1(n_1106_o_0),
    .A2(n_904_o_0),
    .B(n_1109_o_0),
    .C(net14),
    .Y(n_1110_o_0));
 XNOR2xp5_ASAP7_75t_R n_11100 (.A(_01018_),
    .B(n_11099_o_0),
    .Y(n_11100_o_0));
 NOR2xp33_ASAP7_75t_R n_11101 (.A(n_4339_o_0),
    .B(n_11100_o_0),
    .Y(n_11101_o_0));
 NOR2xp33_ASAP7_75t_R n_11102 (.A(_00705_),
    .B(net),
    .Y(n_11102_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11103 (.A1(n_4339_o_0),
    .A2(n_11100_o_0),
    .B(n_11101_o_0),
    .C(net),
    .D(n_11102_o_0),
    .Y(n_11103_o_0));
 NAND2xp33_ASAP7_75t_R n_11104 (.A(_00930_),
    .B(n_11103_o_0),
    .Y(n_11104_o_0));
 OAI21xp33_ASAP7_75t_R n_11105 (.A1(_00930_),
    .A2(n_11103_o_0),
    .B(n_11104_o_0),
    .Y(n_11105_o_0));
 INVx1_ASAP7_75t_R n_11106 (.A(n_11105_o_0),
    .Y(n_11106_o_0));
 XNOR2xp5_ASAP7_75t_R n_11107 (.A(_01057_),
    .B(_01065_),
    .Y(n_11107_o_0));
 XNOR2xp5_ASAP7_75t_R n_11108 (.A(_01103_),
    .B(n_11107_o_0),
    .Y(n_11108_o_0));
 XOR2xp5_ASAP7_75t_R n_11109 (.A(_01016_),
    .B(_01017_),
    .Y(n_11109_o_0));
 INVx1_ASAP7_75t_R n_1111 (.A(n_1012_o_0),
    .Y(n_1111_o_0));
 NOR2xp33_ASAP7_75t_R n_11110 (.A(n_11109_o_0),
    .B(n_11108_o_0),
    .Y(n_11110_o_0));
 NOR2xp33_ASAP7_75t_R n_11111 (.A(_00706_),
    .B(net),
    .Y(n_11111_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11112 (.A1(n_11108_o_0),
    .A2(n_11109_o_0),
    .B(n_11110_o_0),
    .C(net39),
    .D(n_11111_o_0),
    .Y(n_11112_o_0));
 INVx1_ASAP7_75t_R n_11113 (.A(_00929_),
    .Y(n_11113_o_0));
 NAND2xp33_ASAP7_75t_R n_11114 (.A(n_11113_o_0),
    .B(n_11112_o_0),
    .Y(n_11114_o_0));
 OAI21xp5_ASAP7_75t_R n_11115 (.A1(n_11112_o_0),
    .A2(n_11113_o_0),
    .B(n_11114_o_0),
    .Y(n_11115_o_0));
 NAND2xp33_ASAP7_75t_R n_11116 (.A(n_4230_o_0),
    .B(n_4201_o_0),
    .Y(n_11116_o_0));
 OAI21xp33_ASAP7_75t_R n_11117 (.A1(n_4201_o_0),
    .A2(n_4230_o_0),
    .B(n_11116_o_0),
    .Y(n_11117_o_0));
 INVx1_ASAP7_75t_R n_11118 (.A(_01106_),
    .Y(n_11118_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11119 (.A1(n_4230_o_0),
    .A2(n_4201_o_0),
    .B(n_11116_o_0),
    .C(n_11118_o_0),
    .Y(n_11119_o_0));
 OAI21xp33_ASAP7_75t_R n_1112 (.A1(n_907_o_0),
    .A2(n_1111_o_0),
    .B(n_1062_o_0),
    .Y(n_1112_o_0));
 INVx1_ASAP7_75t_R n_11120 (.A(n_11119_o_0),
    .Y(n_11120_o_0));
 OAI21xp33_ASAP7_75t_R n_11121 (.A1(_01106_),
    .A2(n_11117_o_0),
    .B(n_11120_o_0),
    .Y(n_11121_o_0));
 INVx1_ASAP7_75t_R n_11122 (.A(_00638_),
    .Y(n_11122_o_0));
 OAI21xp33_ASAP7_75t_R n_11123 (.A1(net39),
    .A2(n_11122_o_0),
    .B(_00924_),
    .Y(n_11123_o_0));
 NOR2xp33_ASAP7_75t_R n_11124 (.A(_01106_),
    .B(n_11117_o_0),
    .Y(n_11124_o_0));
 AOI21xp33_ASAP7_75t_R n_11125 (.A1(n_11122_o_0),
    .A2(n_3021_o_0),
    .B(_00924_),
    .Y(n_11125_o_0));
 OAI31xp33_ASAP7_75t_R n_11126 (.A1(n_3021_o_0),
    .A2(n_11124_o_0),
    .A3(n_11119_o_0),
    .B(n_11125_o_0),
    .Y(n_11126_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11127 (.A1(n_11121_o_0),
    .A2(net39),
    .B(n_11123_o_0),
    .C(n_11126_o_0),
    .Y(n_11127_o_0));
 XNOR2xp5_ASAP7_75t_R n_11128 (.A(_01061_),
    .B(n_4201_o_0),
    .Y(n_11128_o_0));
 XNOR2xp5_ASAP7_75t_R n_11129 (.A(n_4185_o_0),
    .B(n_8900_o_0),
    .Y(n_11129_o_0));
 OAI21xp33_ASAP7_75t_R n_1113 (.A1(n_989_o_0),
    .A2(n_942_o_0),
    .B(n_903_o_0),
    .Y(n_1113_o_0));
 XNOR2xp5_ASAP7_75t_R n_11130 (.A(n_11128_o_0),
    .B(n_11129_o_0),
    .Y(n_11130_o_0));
 OAI21xp33_ASAP7_75t_R n_11131 (.A1(_00637_),
    .A2(net39),
    .B(_00925_),
    .Y(n_11131_o_0));
 INVx1_ASAP7_75t_R n_11132 (.A(n_11131_o_0),
    .Y(n_11132_o_0));
 AOI21xp33_ASAP7_75t_R n_11133 (.A1(_00637_),
    .A2(net3),
    .B(_00925_),
    .Y(n_11133_o_0));
 INVx1_ASAP7_75t_R n_11134 (.A(n_11133_o_0),
    .Y(n_11134_o_0));
 AOI21xp33_ASAP7_75t_R n_11135 (.A1(net39),
    .A2(n_11130_o_0),
    .B(n_11134_o_0),
    .Y(n_11135_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_11136 (.A1(n_3021_o_0),
    .A2(n_11130_o_0),
    .B(n_11132_o_0),
    .C(n_11135_o_0),
    .Y(n_11136_o_0));
 NOR2xp33_ASAP7_75t_R n_11137 (.A(n_11127_o_0),
    .B(n_11136_o_0),
    .Y(n_11137_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11138 (.A1(_01106_),
    .A2(n_11117_o_0),
    .B(n_11124_o_0),
    .C(net77),
    .D(n_11123_o_0),
    .Y(n_11138_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_11139 (.A1(net5),
    .A2(n_11121_o_0),
    .B(n_11125_o_0),
    .C(n_11138_o_0),
    .Y(n_11139_o_0));
 AO21x1_ASAP7_75t_R n_1114 (.A1(n_887_o_0),
    .A2(n_877_o_0),
    .B(n_1113_o_0),
    .Y(n_1114_o_0));
 INVx1_ASAP7_75t_R n_11140 (.A(_00926_),
    .Y(n_11140_o_0));
 XNOR2xp5_ASAP7_75t_R n_11141 (.A(_01013_),
    .B(_01100_),
    .Y(n_11141_o_0));
 XNOR2xp5_ASAP7_75t_R n_11142 (.A(_01062_),
    .B(n_11141_o_0),
    .Y(n_11142_o_0));
 NAND2xp33_ASAP7_75t_R n_11143 (.A(n_8916_o_0),
    .B(n_11142_o_0),
    .Y(n_11143_o_0));
 OAI21xp33_ASAP7_75t_R n_11144 (.A1(n_8916_o_0),
    .A2(n_11142_o_0),
    .B(n_11143_o_0),
    .Y(n_11144_o_0));
 NOR2xp33_ASAP7_75t_R n_11145 (.A(_00639_),
    .B(net77),
    .Y(n_11145_o_0));
 AOI21xp33_ASAP7_75t_R n_11146 (.A1(net39),
    .A2(n_11144_o_0),
    .B(n_11145_o_0),
    .Y(n_11146_o_0));
 OR2x2_ASAP7_75t_R n_11147 (.A(_01014_),
    .B(_01054_),
    .Y(n_11147_o_0));
 NAND2xp33_ASAP7_75t_R n_11148 (.A(_01014_),
    .B(_01054_),
    .Y(n_11148_o_0));
 AO21x1_ASAP7_75t_R n_11149 (.A1(n_11147_o_0),
    .A2(n_11148_o_0),
    .B(n_11142_o_0),
    .Y(n_11149_o_0));
 OAI211xp5_ASAP7_75t_R n_1115 (.A1(n_903_o_0),
    .A2(n_1112_o_0),
    .B(n_1114_o_0),
    .C(net16),
    .Y(n_1115_o_0));
 INVx1_ASAP7_75t_R n_11150 (.A(n_11145_o_0),
    .Y(n_11150_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11151 (.A1(n_11143_o_0),
    .A2(n_11149_o_0),
    .B(n_3021_o_0),
    .C(n_11150_o_0),
    .D(n_11140_o_0),
    .Y(n_11151_o_0));
 AOI21x1_ASAP7_75t_R n_11152 (.A1(n_11146_o_0),
    .A2(n_11140_o_0),
    .B(n_11151_o_0),
    .Y(n_11152_o_0));
 XNOR2xp5_ASAP7_75t_R n_11153 (.A(_01063_),
    .B(n_4246_o_0),
    .Y(n_11153_o_0));
 XOR2xp5_ASAP7_75t_R n_11154 (.A(n_11153_o_0),
    .B(n_8932_o_0),
    .Y(n_11154_o_0));
 NOR2xp33_ASAP7_75t_R n_11155 (.A(_00708_),
    .B(net39),
    .Y(n_11155_o_0));
 AOI21xp33_ASAP7_75t_R n_11156 (.A1(net39),
    .A2(n_11154_o_0),
    .B(n_11155_o_0),
    .Y(n_11156_o_0));
 XNOR2xp5_ASAP7_75t_R n_11157 (.A(n_11153_o_0),
    .B(n_8932_o_0),
    .Y(n_11157_o_0));
 INVx1_ASAP7_75t_R n_11158 (.A(n_11155_o_0),
    .Y(n_11158_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11159 (.A1(net2),
    .A2(n_11157_o_0),
    .B(n_11158_o_0),
    .C(_00927_),
    .Y(n_11159_o_0));
 NAND3xp33_ASAP7_75t_R n_1116 (.A(n_1110_o_0),
    .B(n_930_o_0),
    .C(n_1115_o_0),
    .Y(n_1116_o_0));
 AO21x1_ASAP7_75t_R n_11160 (.A1(_00927_),
    .A2(n_11156_o_0),
    .B(n_11159_o_0),
    .Y(n_11160_o_0));
 OAI21xp33_ASAP7_75t_R n_11161 (.A1(n_11139_o_0),
    .A2(n_11152_o_0),
    .B(n_11160_o_0),
    .Y(n_11161_o_0));
 AO21x1_ASAP7_75t_R n_11162 (.A1(n_11146_o_0),
    .A2(n_11140_o_0),
    .B(n_11151_o_0),
    .Y(n_11162_o_0));
 INVx1_ASAP7_75t_R n_11163 (.A(_00927_),
    .Y(n_11163_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11164 (.A1(net9),
    .A2(n_11157_o_0),
    .B(n_11158_o_0),
    .C(n_11163_o_0),
    .Y(n_11164_o_0));
 AO21x1_ASAP7_75t_R n_11165 (.A1(n_11163_o_0),
    .A2(n_11156_o_0),
    .B(n_11164_o_0),
    .Y(n_11165_o_0));
 OAI21xp33_ASAP7_75t_R n_11166 (.A1(net58),
    .A2(n_11162_o_0),
    .B(n_11165_o_0),
    .Y(n_11166_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11167 (.A1(n_11121_o_0),
    .A2(net),
    .B(n_11123_o_0),
    .C(n_11126_o_0),
    .Y(n_11167_o_0));
 NAND2xp33_ASAP7_75t_R n_11168 (.A(_01061_),
    .B(n_4213_o_0),
    .Y(n_11168_o_0));
 OAI21xp33_ASAP7_75t_R n_11169 (.A1(_01061_),
    .A2(n_4213_o_0),
    .B(n_11168_o_0),
    .Y(n_11169_o_0));
 OAI311xp33_ASAP7_75t_R n_1117 (.A1(n_930_o_0),
    .A2(n_1099_o_0),
    .A3(n_1105_o_0),
    .B1(n_1116_o_0),
    .C1(n_972_o_0),
    .Y(n_1117_o_0));
 XNOR2xp5_ASAP7_75t_R n_11170 (.A(n_11129_o_0),
    .B(n_11169_o_0),
    .Y(n_11170_o_0));
 AOI21xp33_ASAP7_75t_R n_11171 (.A1(net),
    .A2(n_11170_o_0),
    .B(n_11131_o_0),
    .Y(n_11171_o_0));
 NOR3xp33_ASAP7_75t_R n_11172 (.A(n_11167_o_0),
    .B(n_11171_o_0),
    .C(n_11135_o_0),
    .Y(n_11172_o_0));
 XNOR2xp5_ASAP7_75t_R n_11173 (.A(_01064_),
    .B(n_4268_o_0),
    .Y(n_11173_o_0));
 NOR2xp33_ASAP7_75t_R n_11174 (.A(n_11173_o_0),
    .B(n_8882_o_0),
    .Y(n_11174_o_0));
 NOR2xp33_ASAP7_75t_R n_11175 (.A(_00707_),
    .B(net39),
    .Y(n_11175_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11176 (.A1(n_8882_o_0),
    .A2(n_11173_o_0),
    .B(n_11174_o_0),
    .C(net77),
    .D(n_11175_o_0),
    .Y(n_11176_o_0));
 HAxp5_ASAP7_75t_R n_11177 (.A(n_11176_o_0),
    .B(n_1883_o_0),
    .CON(n_11177_o_0),
    .SN(n_11177_o_1));
 OA21x2_ASAP7_75t_R n_11178 (.A1(n_11166_o_0),
    .A2(n_11172_o_0),
    .B(n_11177_o_1),
    .Y(n_11178_o_0));
 NAND3xp33_ASAP7_75t_R n_11179 (.A(n_11136_o_0),
    .B(n_11152_o_0),
    .C(n_11127_o_0),
    .Y(n_11179_o_0));
 OAI31xp33_ASAP7_75t_R n_1118 (.A1(n_972_o_0),
    .A2(n_1078_o_0),
    .A3(n_1092_o_0),
    .B(n_1117_o_0),
    .Y(n_1118_o_0));
 OAI21xp33_ASAP7_75t_R n_11180 (.A1(net9),
    .A2(n_11170_o_0),
    .B(n_11133_o_0),
    .Y(n_11180_o_0));
 OAI21xp33_ASAP7_75t_R n_11181 (.A1(net9),
    .A2(n_11130_o_0),
    .B(n_11132_o_0),
    .Y(n_11181_o_0));
 AOI21xp33_ASAP7_75t_R n_11182 (.A1(n_11180_o_0),
    .A2(n_11181_o_0),
    .B(n_11127_o_0),
    .Y(n_11182_o_0));
 INVx1_ASAP7_75t_R n_11183 (.A(n_11138_o_0),
    .Y(n_11183_o_0));
 AOI211xp5_ASAP7_75t_R n_11184 (.A1(n_11183_o_0),
    .A2(n_11126_o_0),
    .B(n_11171_o_0),
    .C(n_11135_o_0),
    .Y(n_11184_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11185 (.A1(n_11182_o_0),
    .A2(n_11184_o_0),
    .B(n_11162_o_0),
    .C(n_11165_o_0),
    .Y(n_11185_o_0));
 OAI21xp33_ASAP7_75t_R n_11186 (.A1(n_11135_o_0),
    .A2(n_11171_o_0),
    .B(n_11127_o_0),
    .Y(n_11186_o_0));
 INVx1_ASAP7_75t_R n_11187 (.A(n_11186_o_0),
    .Y(n_11187_o_0));
 OAI21xp33_ASAP7_75t_R n_11188 (.A1(n_11135_o_0),
    .A2(n_11171_o_0),
    .B(n_11139_o_0),
    .Y(n_11188_o_0));
 NOR2xp33_ASAP7_75t_R n_11189 (.A(n_11188_o_0),
    .B(n_11162_o_0),
    .Y(n_11189_o_0));
 INVx1_ASAP7_75t_R n_1119 (.A(n_909_o_0),
    .Y(n_1119_o_0));
 AOI21x1_ASAP7_75t_R n_11190 (.A1(n_11163_o_0),
    .A2(n_11156_o_0),
    .B(n_11164_o_0),
    .Y(n_11190_o_0));
 AOI211xp5_ASAP7_75t_R n_11191 (.A1(n_11162_o_0),
    .A2(n_11187_o_0),
    .B(n_11189_o_0),
    .C(n_11190_o_0),
    .Y(n_11191_o_0));
 OAI21xp33_ASAP7_75t_R n_11192 (.A1(n_11176_o_0),
    .A2(n_1883_o_0),
    .B(n_11177_o_0),
    .Y(n_11192_o_0));
 AOI211xp5_ASAP7_75t_R n_11193 (.A1(n_11179_o_0),
    .A2(n_11185_o_0),
    .B(n_11191_o_0),
    .C(n_11192_o_0),
    .Y(n_11193_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11194 (.A1(n_11137_o_0),
    .A2(n_11161_o_0),
    .B(n_11178_o_0),
    .C(n_11193_o_0),
    .Y(n_11194_o_0));
 INVx1_ASAP7_75t_R n_11195 (.A(n_11189_o_0),
    .Y(n_11195_o_0));
 NAND3xp33_ASAP7_75t_R n_11196 (.A(n_11127_o_0),
    .B(n_11180_o_0),
    .C(n_11181_o_0),
    .Y(n_11196_o_0));
 OAI21xp5_ASAP7_75t_R n_11197 (.A1(n_11136_o_0),
    .A2(n_11127_o_0),
    .B(n_11196_o_0),
    .Y(n_11197_o_0));
 AOI21xp33_ASAP7_75t_R n_11198 (.A1(n_11162_o_0),
    .A2(n_11197_o_0),
    .B(n_11190_o_0),
    .Y(n_11198_o_0));
 AOI211xp5_ASAP7_75t_R n_11199 (.A1(n_11154_o_0),
    .A2(net),
    .B(n_11163_o_0),
    .C(n_11155_o_0),
    .Y(n_11199_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1120 (.A1(n_1119_o_0),
    .A2(n_994_o_0),
    .B(n_877_o_0),
    .C(n_829_o_0),
    .Y(n_1120_o_0));
 NOR2xp33_ASAP7_75t_R n_11200 (.A(n_11159_o_0),
    .B(n_11199_o_0),
    .Y(n_11200_o_0));
 NAND2xp33_ASAP7_75t_R n_11201 (.A(n_11188_o_0),
    .B(n_11162_o_0),
    .Y(n_11201_o_0));
 INVx1_ASAP7_75t_R n_11202 (.A(n_11192_o_0),
    .Y(n_11202_o_0));
 OAI21xp33_ASAP7_75t_R n_11203 (.A1(n_11200_o_0),
    .A2(n_11201_o_0),
    .B(n_11202_o_0),
    .Y(n_11203_o_0));
 AOI21xp33_ASAP7_75t_R n_11204 (.A1(n_11195_o_0),
    .A2(n_11198_o_0),
    .B(n_11203_o_0),
    .Y(n_11204_o_0));
 NAND3xp33_ASAP7_75t_R n_11205 (.A(n_11160_o_0),
    .B(n_11186_o_0),
    .C(net65),
    .Y(n_11205_o_0));
 NAND2xp33_ASAP7_75t_R n_11206 (.A(n_11152_o_0),
    .B(n_11136_o_0),
    .Y(n_11206_o_0));
 INVx1_ASAP7_75t_R n_11207 (.A(n_11182_o_0),
    .Y(n_11207_o_0));
 AOI31xp33_ASAP7_75t_R n_11208 (.A1(n_11162_o_0),
    .A2(n_11207_o_0),
    .A3(n_11196_o_0),
    .B(n_11200_o_0),
    .Y(n_11208_o_0));
 AOI21xp33_ASAP7_75t_R n_11209 (.A1(n_11152_o_0),
    .A2(n_11197_o_0),
    .B(n_11190_o_0),
    .Y(n_11209_o_0));
 NOR2xp33_ASAP7_75t_R n_1121 (.A(n_877_o_0),
    .B(n_938_o_0),
    .Y(n_1121_o_0));
 AOI21xp33_ASAP7_75t_R n_11210 (.A1(n_11206_o_0),
    .A2(n_11208_o_0),
    .B(n_11209_o_0),
    .Y(n_11210_o_0));
 NAND2xp33_ASAP7_75t_R n_11211 (.A(_00929_),
    .B(n_11112_o_0),
    .Y(n_11211_o_0));
 OAI21xp33_ASAP7_75t_R n_11212 (.A1(_00929_),
    .A2(n_11112_o_0),
    .B(n_11211_o_0),
    .Y(n_11212_o_0));
 OAI21xp33_ASAP7_75t_R n_11213 (.A1(n_11202_o_0),
    .A2(n_11210_o_0),
    .B(n_11212_o_0),
    .Y(n_11213_o_0));
 AOI21xp33_ASAP7_75t_R n_11214 (.A1(n_11204_o_0),
    .A2(n_11205_o_0),
    .B(n_11213_o_0),
    .Y(n_11214_o_0));
 XOR2xp5_ASAP7_75t_R n_11215 (.A(_01018_),
    .B(_01105_),
    .Y(n_11215_o_0));
 XNOR2xp5_ASAP7_75t_R n_11216 (.A(_01019_),
    .B(n_11215_o_0),
    .Y(n_11216_o_0));
 NOR2xp33_ASAP7_75t_R n_11217 (.A(n_4395_o_0),
    .B(n_11216_o_0),
    .Y(n_11217_o_0));
 NOR2xp33_ASAP7_75t_R n_11218 (.A(_00704_),
    .B(net),
    .Y(n_11218_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11219 (.A1(n_4395_o_0),
    .A2(n_11216_o_0),
    .B(n_11217_o_0),
    .C(net),
    .D(n_11218_o_0),
    .Y(n_11219_o_0));
 OAI21xp33_ASAP7_75t_R n_1122 (.A1(n_1006_o_0),
    .A2(n_890_o_0),
    .B(net16),
    .Y(n_1122_o_0));
 XNOR2xp5_ASAP7_75t_R n_11220 (.A(_00931_),
    .B(n_11219_o_0),
    .Y(n_11220_o_0));
 INVx1_ASAP7_75t_R n_11221 (.A(n_11220_o_0),
    .Y(n_11221_o_0));
 AOI211xp5_ASAP7_75t_R n_11222 (.A1(n_11115_o_0),
    .A2(n_11194_o_0),
    .B(n_11214_o_0),
    .C(n_11221_o_0),
    .Y(n_11222_o_0));
 INVx1_ASAP7_75t_R n_11223 (.A(n_11212_o_0),
    .Y(n_11223_o_0));
 INVx1_ASAP7_75t_R n_11224 (.A(n_11177_o_1),
    .Y(n_11224_o_0));
 NOR3xp33_ASAP7_75t_R n_11225 (.A(n_11165_o_0),
    .B(n_11188_o_0),
    .C(net65),
    .Y(n_11225_o_0));
 INVx1_ASAP7_75t_R n_11226 (.A(n_11225_o_0),
    .Y(n_11226_o_0));
 AOI31xp33_ASAP7_75t_R n_11227 (.A1(net58),
    .A2(net35),
    .A3(n_11162_o_0),
    .B(n_11160_o_0),
    .Y(n_11227_o_0));
 OAI21xp33_ASAP7_75t_R n_11228 (.A1(n_11162_o_0),
    .A2(n_11187_o_0),
    .B(n_11227_o_0),
    .Y(n_11228_o_0));
 NOR4xp25_ASAP7_75t_R n_11229 (.A(n_11152_o_0),
    .B(n_11167_o_0),
    .C(n_11135_o_0),
    .D(n_11171_o_0),
    .Y(n_11229_o_0));
 AOI21xp33_ASAP7_75t_R n_1123 (.A1(n_1121_o_0),
    .A2(n_953_o_0),
    .B(n_1122_o_0),
    .Y(n_1123_o_0));
 OAI21xp33_ASAP7_75t_R n_11230 (.A1(n_11162_o_0),
    .A2(n_11186_o_0),
    .B(n_11160_o_0),
    .Y(n_11230_o_0));
 NAND2xp33_ASAP7_75t_R n_11231 (.A(n_11200_o_0),
    .B(n_11162_o_0),
    .Y(n_11231_o_0));
 OAI221xp5_ASAP7_75t_R n_11232 (.A1(n_11229_o_0),
    .A2(n_11230_o_0),
    .B1(n_11231_o_0),
    .B2(n_11188_o_0),
    .C(n_11192_o_0),
    .Y(n_11232_o_0));
 INVx1_ASAP7_75t_R n_11233 (.A(n_11232_o_0),
    .Y(n_11233_o_0));
 AOI31xp33_ASAP7_75t_R n_11234 (.A1(n_11224_o_0),
    .A2(n_11226_o_0),
    .A3(n_11228_o_0),
    .B(n_11233_o_0),
    .Y(n_11234_o_0));
 AOI21xp33_ASAP7_75t_R n_11235 (.A1(n_11139_o_0),
    .A2(n_11136_o_0),
    .B(n_11162_o_0),
    .Y(n_11235_o_0));
 NOR3xp33_ASAP7_75t_R n_11236 (.A(n_11229_o_0),
    .B(n_11235_o_0),
    .C(n_11165_o_0),
    .Y(n_11236_o_0));
 NAND2xp33_ASAP7_75t_R n_11237 (.A(n_11152_o_0),
    .B(n_11190_o_0),
    .Y(n_11237_o_0));
 NOR2xp33_ASAP7_75t_R n_11238 (.A(n_11188_o_0),
    .B(n_11237_o_0),
    .Y(n_11238_o_0));
 NAND2xp33_ASAP7_75t_R n_11239 (.A(n_11127_o_0),
    .B(n_11152_o_0),
    .Y(n_11239_o_0));
 AOI21xp33_ASAP7_75t_R n_1124 (.A1(n_942_o_0),
    .A2(n_1120_o_0),
    .B(n_1123_o_0),
    .Y(n_1124_o_0));
 NAND2xp33_ASAP7_75t_R n_11240 (.A(n_11188_o_0),
    .B(n_11162_o_0),
    .Y(n_11240_o_0));
 AOI21xp33_ASAP7_75t_R n_11241 (.A1(n_11239_o_0),
    .A2(n_11240_o_0),
    .B(n_11160_o_0),
    .Y(n_11241_o_0));
 NOR4xp25_ASAP7_75t_R n_11242 (.A(n_11236_o_0),
    .B(n_11238_o_0),
    .C(n_11241_o_0),
    .D(net49),
    .Y(n_11242_o_0));
 OAI211xp5_ASAP7_75t_R n_11243 (.A1(n_11136_o_0),
    .A2(net68),
    .B(n_11196_o_0),
    .C(n_11152_o_0),
    .Y(n_11243_o_0));
 INVx1_ASAP7_75t_R n_11244 (.A(n_11243_o_0),
    .Y(n_11244_o_0));
 NAND2xp33_ASAP7_75t_R n_11245 (.A(net35),
    .B(n_11162_o_0),
    .Y(n_11245_o_0));
 OAI21xp33_ASAP7_75t_R n_11246 (.A1(n_11160_o_0),
    .A2(n_11245_o_0),
    .B(n_11192_o_0),
    .Y(n_11246_o_0));
 AOI21xp33_ASAP7_75t_R n_11247 (.A1(n_11190_o_0),
    .A2(n_11244_o_0),
    .B(n_11246_o_0),
    .Y(n_11247_o_0));
 OAI31xp33_ASAP7_75t_R n_11248 (.A1(n_11115_o_0),
    .A2(n_11242_o_0),
    .A3(n_11247_o_0),
    .B(n_11221_o_0),
    .Y(n_11248_o_0));
 AOI21xp33_ASAP7_75t_R n_11249 (.A1(n_11223_o_0),
    .A2(n_11234_o_0),
    .B(n_11248_o_0),
    .Y(n_11249_o_0));
 OAI21xp33_ASAP7_75t_R n_1125 (.A1(n_881_o_0),
    .A2(n_1044_o_0),
    .B(n_1051_o_0),
    .Y(n_1125_o_0));
 NAND2xp5_ASAP7_75t_R n_11250 (.A(n_11181_o_0),
    .B(n_11180_o_0),
    .Y(n_11250_o_0));
 AOI21xp33_ASAP7_75t_R n_11251 (.A1(n_11139_o_0),
    .A2(n_11250_o_0),
    .B(n_11162_o_0),
    .Y(n_11251_o_0));
 INVx1_ASAP7_75t_R n_11252 (.A(n_11251_o_0),
    .Y(n_11252_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11253 (.A1(n_11188_o_0),
    .A2(net65),
    .B(n_11252_o_0),
    .C(n_11165_o_0),
    .Y(n_11253_o_0));
 INVx1_ASAP7_75t_R n_11254 (.A(n_11253_o_0),
    .Y(n_11254_o_0));
 OAI21xp33_ASAP7_75t_R n_11255 (.A1(net37),
    .A2(n_11250_o_0),
    .B(n_11162_o_0),
    .Y(n_11255_o_0));
 AOI21xp33_ASAP7_75t_R n_11256 (.A1(n_11165_o_0),
    .A2(n_11255_o_0),
    .B(n_11224_o_0),
    .Y(n_11256_o_0));
 NOR2xp33_ASAP7_75t_R n_11257 (.A(n_11186_o_0),
    .B(n_11162_o_0),
    .Y(n_11257_o_0));
 INVx1_ASAP7_75t_R n_11258 (.A(n_11257_o_0),
    .Y(n_11258_o_0));
 AOI21xp33_ASAP7_75t_R n_11259 (.A1(n_11139_o_0),
    .A2(n_11162_o_0),
    .B(n_11190_o_0),
    .Y(n_11259_o_0));
 OAI31xp33_ASAP7_75t_R n_1126 (.A1(net32),
    .A2(n_917_o_0),
    .A3(n_877_o_0),
    .B(n_1125_o_0),
    .Y(n_1126_o_0));
 OAI21xp33_ASAP7_75t_R n_11260 (.A1(n_11152_o_0),
    .A2(n_11250_o_0),
    .B(n_11160_o_0),
    .Y(n_11260_o_0));
 OAI21xp33_ASAP7_75t_R n_11261 (.A1(n_11260_o_0),
    .A2(n_11244_o_0),
    .B(n_11202_o_0),
    .Y(n_11261_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11262 (.A1(n_11258_o_0),
    .A2(n_11259_o_0),
    .B(n_11261_o_0),
    .C(n_11115_o_0),
    .Y(n_11262_o_0));
 AOI21xp33_ASAP7_75t_R n_11263 (.A1(n_11162_o_0),
    .A2(n_11197_o_0),
    .B(n_11160_o_0),
    .Y(n_11263_o_0));
 NAND2xp33_ASAP7_75t_R n_11264 (.A(n_11139_o_0),
    .B(n_11136_o_0),
    .Y(n_11264_o_0));
 OAI32xp33_ASAP7_75t_R n_11265 (.A1(n_11165_o_0),
    .A2(n_11186_o_0),
    .A3(n_11152_o_0),
    .B1(n_11237_o_0),
    .B2(n_11264_o_0),
    .Y(n_11265_o_0));
 INVx1_ASAP7_75t_R n_11266 (.A(n_11115_o_0),
    .Y(n_11266_o_0));
 NAND4xp25_ASAP7_75t_R n_11267 (.A(n_11190_o_0),
    .B(n_11152_o_0),
    .C(n_11136_o_0),
    .D(n_11139_o_0),
    .Y(n_11267_o_0));
 NAND3xp33_ASAP7_75t_R n_11268 (.A(n_11162_o_0),
    .B(net68),
    .C(n_11136_o_0),
    .Y(n_11268_o_0));
 AOI21xp33_ASAP7_75t_R n_11269 (.A1(n_11139_o_0),
    .A2(n_11152_o_0),
    .B(n_11160_o_0),
    .Y(n_11269_o_0));
 AOI311xp33_ASAP7_75t_R n_1127 (.A1(n_877_o_0),
    .A2(n_882_o_0),
    .A3(n_865_o_0),
    .B(n_891_o_0),
    .C(n_911_o_0),
    .Y(n_1127_o_0));
 AOI21xp33_ASAP7_75t_R n_11270 (.A1(n_11268_o_0),
    .A2(n_11269_o_0),
    .B(n_11177_o_1),
    .Y(n_11270_o_0));
 NAND2xp33_ASAP7_75t_R n_11271 (.A(n_11267_o_0),
    .B(n_11270_o_0),
    .Y(n_11271_o_0));
 OAI311xp33_ASAP7_75t_R n_11272 (.A1(n_11202_o_0),
    .A2(n_11263_o_0),
    .A3(n_11265_o_0),
    .B1(n_11266_o_0),
    .C1(n_11271_o_0),
    .Y(n_11272_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11273 (.A1(n_11254_o_0),
    .A2(n_11256_o_0),
    .B(n_11262_o_0),
    .C(n_11272_o_0),
    .Y(n_11273_o_0));
 OAI21xp33_ASAP7_75t_R n_11274 (.A1(n_11152_o_0),
    .A2(net68),
    .B(n_11160_o_0),
    .Y(n_11274_o_0));
 AOI21xp33_ASAP7_75t_R n_11275 (.A1(net65),
    .A2(n_11172_o_0),
    .B(n_11274_o_0),
    .Y(n_11275_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11276 (.A1(n_11207_o_0),
    .A2(n_11196_o_0),
    .B(n_11152_o_0),
    .C(n_11165_o_0),
    .Y(n_11276_o_0));
 NOR2xp33_ASAP7_75t_R n_11277 (.A(n_11139_o_0),
    .B(n_11250_o_0),
    .Y(n_11277_o_0));
 NOR2xp33_ASAP7_75t_R n_11278 (.A(n_11162_o_0),
    .B(n_11277_o_0),
    .Y(n_11278_o_0));
 OAI21xp33_ASAP7_75t_R n_11279 (.A1(n_11276_o_0),
    .A2(n_11278_o_0),
    .B(net49),
    .Y(n_11279_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1128 (.A1(n_1126_o_0),
    .A2(n_1030_o_0),
    .B(net15),
    .C(n_1127_o_0),
    .Y(n_1128_o_0));
 AOI21xp33_ASAP7_75t_R n_11280 (.A1(net58),
    .A2(n_11152_o_0),
    .B(n_11200_o_0),
    .Y(n_11280_o_0));
 INVx1_ASAP7_75t_R n_11281 (.A(n_11280_o_0),
    .Y(n_11281_o_0));
 NAND4xp25_ASAP7_75t_R n_11282 (.A(n_11183_o_0),
    .B(n_11180_o_0),
    .C(n_11181_o_0),
    .D(n_11126_o_0),
    .Y(n_11282_o_0));
 OAI211xp5_ASAP7_75t_R n_11283 (.A1(n_11162_o_0),
    .A2(n_11282_o_0),
    .B(n_11255_o_0),
    .C(n_11165_o_0),
    .Y(n_11283_o_0));
 AOI31xp33_ASAP7_75t_R n_11284 (.A1(n_11281_o_0),
    .A2(n_11283_o_0),
    .A3(n_11202_o_0),
    .B(n_11266_o_0),
    .Y(n_11284_o_0));
 OAI21xp33_ASAP7_75t_R n_11285 (.A1(n_11275_o_0),
    .A2(n_11279_o_0),
    .B(n_11284_o_0),
    .Y(n_11285_o_0));
 AOI211xp5_ASAP7_75t_R n_11286 (.A1(n_11162_o_0),
    .A2(net37),
    .B(n_11165_o_0),
    .C(net35),
    .Y(n_11286_o_0));
 INVx1_ASAP7_75t_R n_11287 (.A(n_11286_o_0),
    .Y(n_11287_o_0));
 AOI21xp33_ASAP7_75t_R n_11288 (.A1(n_11287_o_0),
    .A2(n_11270_o_0),
    .B(n_11115_o_0),
    .Y(n_11288_o_0));
 AOI21xp33_ASAP7_75t_R n_11289 (.A1(n_11152_o_0),
    .A2(n_11172_o_0),
    .B(n_11200_o_0),
    .Y(n_11289_o_0));
 AOI21xp33_ASAP7_75t_R n_1129 (.A1(n_904_o_0),
    .A2(n_1128_o_0),
    .B(n_930_o_0),
    .Y(n_1129_o_0));
 INVx1_ASAP7_75t_R n_11290 (.A(n_11289_o_0),
    .Y(n_11290_o_0));
 NAND2xp33_ASAP7_75t_R n_11291 (.A(n_11127_o_0),
    .B(n_11136_o_0),
    .Y(n_11291_o_0));
 NAND2xp33_ASAP7_75t_R n_11292 (.A(n_11162_o_0),
    .B(n_11291_o_0),
    .Y(n_11292_o_0));
 AOI21xp33_ASAP7_75t_R n_11293 (.A1(n_11269_o_0),
    .A2(n_11292_o_0),
    .B(n_11202_o_0),
    .Y(n_11293_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11294 (.A1(n_11250_o_0),
    .A2(n_11162_o_0),
    .B(n_11290_o_0),
    .C(n_11293_o_0),
    .Y(n_11294_o_0));
 AOI21xp33_ASAP7_75t_R n_11295 (.A1(n_11288_o_0),
    .A2(n_11294_o_0),
    .B(n_11221_o_0),
    .Y(n_11295_o_0));
 XNOR2xp5_ASAP7_75t_R n_11296 (.A(_00930_),
    .B(n_11103_o_0),
    .Y(n_11296_o_0));
 AOI21xp33_ASAP7_75t_R n_11297 (.A1(n_11285_o_0),
    .A2(n_11295_o_0),
    .B(n_11296_o_0),
    .Y(n_11297_o_0));
 OAI21xp33_ASAP7_75t_R n_11298 (.A1(n_11220_o_0),
    .A2(n_11273_o_0),
    .B(n_11297_o_0),
    .Y(n_11298_o_0));
 OAI31xp33_ASAP7_75t_R n_11299 (.A1(n_11106_o_0),
    .A2(n_11222_o_0),
    .A3(n_11249_o_0),
    .B(n_11298_o_0),
    .Y(n_11299_o_0));
 OAI21xp33_ASAP7_75t_R n_1130 (.A1(n_1124_o_0),
    .A2(n_904_o_0),
    .B(n_1129_o_0),
    .Y(n_1130_o_0));
 AOI21xp33_ASAP7_75t_R n_11300 (.A1(n_11165_o_0),
    .A2(n_11206_o_0),
    .B(n_11224_o_0),
    .Y(n_11300_o_0));
 OA21x2_ASAP7_75t_R n_11301 (.A1(net35),
    .A2(net65),
    .B(n_11267_o_0),
    .Y(n_11301_o_0));
 AOI21xp33_ASAP7_75t_R n_11302 (.A1(net65),
    .A2(n_11197_o_0),
    .B(n_11160_o_0),
    .Y(n_11302_o_0));
 AOI211xp5_ASAP7_75t_R n_11303 (.A1(n_11292_o_0),
    .A2(n_11302_o_0),
    .B(n_11236_o_0),
    .C(net49),
    .Y(n_11303_o_0));
 AOI211xp5_ASAP7_75t_R n_11304 (.A1(n_11300_o_0),
    .A2(n_11301_o_0),
    .B(n_11303_o_0),
    .C(n_11106_o_0),
    .Y(n_11304_o_0));
 NOR2xp33_ASAP7_75t_R n_11305 (.A(n_11162_o_0),
    .B(n_11264_o_0),
    .Y(n_11305_o_0));
 AOI21xp33_ASAP7_75t_R n_11306 (.A1(net37),
    .A2(n_11152_o_0),
    .B(n_11200_o_0),
    .Y(n_11306_o_0));
 AOI21xp33_ASAP7_75t_R n_11307 (.A1(n_11306_o_0),
    .A2(n_11240_o_0),
    .B(n_11224_o_0),
    .Y(n_11307_o_0));
 OAI21xp33_ASAP7_75t_R n_11308 (.A1(n_11305_o_0),
    .A2(n_11276_o_0),
    .B(n_11307_o_0),
    .Y(n_11308_o_0));
 NAND2xp33_ASAP7_75t_R n_11309 (.A(net68),
    .B(n_11136_o_0),
    .Y(n_11309_o_0));
 NOR2xp33_ASAP7_75t_R n_1131 (.A(n_1060_o_0),
    .B(n_890_o_0),
    .Y(n_1131_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11310 (.A1(n_11197_o_0),
    .A2(net65),
    .B(n_11161_o_0),
    .C(n_11202_o_0),
    .Y(n_11310_o_0));
 AO21x1_ASAP7_75t_R n_11311 (.A1(n_11259_o_0),
    .A2(n_11309_o_0),
    .B(n_11310_o_0),
    .Y(n_11311_o_0));
 AOI21xp33_ASAP7_75t_R n_11312 (.A1(n_11308_o_0),
    .A2(n_11311_o_0),
    .B(n_11105_o_0),
    .Y(n_11312_o_0));
 NOR3xp33_ASAP7_75t_R n_11313 (.A(n_11304_o_0),
    .B(n_11312_o_0),
    .C(n_11115_o_0),
    .Y(n_11313_o_0));
 NOR2xp33_ASAP7_75t_R n_11314 (.A(n_11152_o_0),
    .B(n_11136_o_0),
    .Y(n_11314_o_0));
 NAND3xp33_ASAP7_75t_R n_11315 (.A(n_11309_o_0),
    .B(n_11160_o_0),
    .C(n_11162_o_0),
    .Y(n_11315_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11316 (.A1(n_11190_o_0),
    .A2(n_11314_o_0),
    .B(n_11315_o_0),
    .C(n_11278_o_0),
    .Y(n_11316_o_0));
 NAND3xp33_ASAP7_75t_R n_11317 (.A(n_11190_o_0),
    .B(net35),
    .C(net58),
    .Y(n_11317_o_0));
 OAI211xp5_ASAP7_75t_R n_11318 (.A1(net37),
    .A2(net35),
    .B(n_11196_o_0),
    .C(n_11162_o_0),
    .Y(n_11318_o_0));
 AOI31xp33_ASAP7_75t_R n_11319 (.A1(net35),
    .A2(net65),
    .A3(net37),
    .B(n_11160_o_0),
    .Y(n_11319_o_0));
 AOI31xp33_ASAP7_75t_R n_1132 (.A1(n_950_o_0),
    .A2(n_1029_o_0),
    .A3(n_878_o_0),
    .B(n_1131_o_0),
    .Y(n_1132_o_0));
 AOI21xp33_ASAP7_75t_R n_11320 (.A1(n_11318_o_0),
    .A2(n_11319_o_0),
    .B(n_11192_o_0),
    .Y(n_11320_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11321 (.A1(n_11317_o_0),
    .A2(net65),
    .B(n_11320_o_0),
    .C(n_11296_o_0),
    .Y(n_11321_o_0));
 OA21x2_ASAP7_75t_R n_11322 (.A1(n_11224_o_0),
    .A2(n_11316_o_0),
    .B(n_11321_o_0),
    .Y(n_11322_o_0));
 INVx1_ASAP7_75t_R n_11323 (.A(n_11137_o_0),
    .Y(n_11323_o_0));
 NAND2xp33_ASAP7_75t_R n_11324 (.A(n_11136_o_0),
    .B(n_11162_o_0),
    .Y(n_11324_o_0));
 NOR3xp33_ASAP7_75t_R n_11325 (.A(n_11172_o_0),
    .B(n_11162_o_0),
    .C(n_11190_o_0),
    .Y(n_11325_o_0));
 AOI31xp33_ASAP7_75t_R n_11326 (.A1(n_11160_o_0),
    .A2(n_11323_o_0),
    .A3(n_11324_o_0),
    .B(n_11325_o_0),
    .Y(n_11326_o_0));
 AO211x2_ASAP7_75t_R n_11327 (.A1(n_11146_o_0),
    .A2(n_11140_o_0),
    .B(n_11151_o_0),
    .C(net68),
    .Y(n_11327_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11328 (.A1(n_11136_o_0),
    .A2(n_11139_o_0),
    .B(n_11152_o_0),
    .C(n_11190_o_0),
    .Y(n_11328_o_0));
 INVx1_ASAP7_75t_R n_11329 (.A(n_11239_o_0),
    .Y(n_11329_o_0));
 OAI21xp33_ASAP7_75t_R n_1133 (.A1(net16),
    .A2(n_1132_o_0),
    .B(n_904_o_0),
    .Y(n_1133_o_0));
 OAI21xp33_ASAP7_75t_R n_11330 (.A1(n_11328_o_0),
    .A2(n_11329_o_0),
    .B(n_11177_o_1),
    .Y(n_11330_o_0));
 AOI21xp33_ASAP7_75t_R n_11331 (.A1(n_11198_o_0),
    .A2(n_11327_o_0),
    .B(n_11330_o_0),
    .Y(n_11331_o_0));
 AOI211xp5_ASAP7_75t_R n_11332 (.A1(n_11202_o_0),
    .A2(n_11326_o_0),
    .B(n_11331_o_0),
    .C(n_11106_o_0),
    .Y(n_11332_o_0));
 NOR3xp33_ASAP7_75t_R n_11333 (.A(n_11322_o_0),
    .B(n_11332_o_0),
    .C(n_11212_o_0),
    .Y(n_11333_o_0));
 OAI21xp33_ASAP7_75t_R n_11334 (.A1(n_11152_o_0),
    .A2(n_11277_o_0),
    .B(n_11190_o_0),
    .Y(n_11334_o_0));
 OAI21xp33_ASAP7_75t_R n_11335 (.A1(n_11251_o_0),
    .A2(n_11334_o_0),
    .B(n_11266_o_0),
    .Y(n_11335_o_0));
 AOI21xp33_ASAP7_75t_R n_11336 (.A1(n_11319_o_0),
    .A2(n_11318_o_0),
    .B(n_11335_o_0),
    .Y(n_11336_o_0));
 NAND2xp33_ASAP7_75t_R n_11337 (.A(n_11165_o_0),
    .B(n_11243_o_0),
    .Y(n_11337_o_0));
 INVx1_ASAP7_75t_R n_11338 (.A(n_11306_o_0),
    .Y(n_11338_o_0));
 OAI21xp33_ASAP7_75t_R n_11339 (.A1(n_11160_o_0),
    .A2(n_11240_o_0),
    .B(n_11115_o_0),
    .Y(n_11339_o_0));
 AOI211xp5_ASAP7_75t_R n_1134 (.A1(n_881_o_0),
    .A2(n_918_o_0),
    .B(n_994_o_0),
    .C(n_878_o_0),
    .Y(n_1134_o_0));
 AOI211xp5_ASAP7_75t_R n_11340 (.A1(n_11337_o_0),
    .A2(n_11338_o_0),
    .B(n_11225_o_0),
    .C(n_11339_o_0),
    .Y(n_11340_o_0));
 INVx1_ASAP7_75t_R n_11341 (.A(n_11206_o_0),
    .Y(n_11341_o_0));
 OAI21xp33_ASAP7_75t_R n_11342 (.A1(n_11161_o_0),
    .A2(n_11341_o_0),
    .B(n_11266_o_0),
    .Y(n_11342_o_0));
 OAI211xp5_ASAP7_75t_R n_11343 (.A1(n_11139_o_0),
    .A2(n_11152_o_0),
    .B(n_11165_o_0),
    .C(net35),
    .Y(n_11343_o_0));
 INVx1_ASAP7_75t_R n_11344 (.A(n_11343_o_0),
    .Y(n_11344_o_0));
 NAND3xp33_ASAP7_75t_R n_11345 (.A(n_11162_o_0),
    .B(net68),
    .C(n_11136_o_0),
    .Y(n_11345_o_0));
 AOI21xp33_ASAP7_75t_R n_11346 (.A1(n_11152_o_0),
    .A2(n_11172_o_0),
    .B(n_11190_o_0),
    .Y(n_11346_o_0));
 AOI21xp33_ASAP7_75t_R n_11347 (.A1(n_11345_o_0),
    .A2(n_11346_o_0),
    .B(n_11212_o_0),
    .Y(n_11347_o_0));
 OAI21xp33_ASAP7_75t_R n_11348 (.A1(n_11189_o_0),
    .A2(n_11274_o_0),
    .B(n_11347_o_0),
    .Y(n_11348_o_0));
 OAI211xp5_ASAP7_75t_R n_11349 (.A1(n_11342_o_0),
    .A2(n_11344_o_0),
    .B(n_11348_o_0),
    .C(n_11105_o_0),
    .Y(n_11349_o_0));
 AOI211xp5_ASAP7_75t_R n_1135 (.A1(n_1107_o_0),
    .A2(n_893_o_0),
    .B(net15),
    .C(n_1134_o_0),
    .Y(n_1135_o_0));
 OAI31xp33_ASAP7_75t_R n_11350 (.A1(n_11105_o_0),
    .A2(n_11336_o_0),
    .A3(n_11340_o_0),
    .B(n_11349_o_0),
    .Y(n_11350_o_0));
 NOR2xp33_ASAP7_75t_R n_11351 (.A(n_11136_o_0),
    .B(n_11162_o_0),
    .Y(n_11351_o_0));
 NOR2xp33_ASAP7_75t_R n_11352 (.A(n_11139_o_0),
    .B(n_11152_o_0),
    .Y(n_11352_o_0));
 INVx1_ASAP7_75t_R n_11353 (.A(n_11352_o_0),
    .Y(n_11353_o_0));
 INVx1_ASAP7_75t_R n_11354 (.A(n_11230_o_0),
    .Y(n_11354_o_0));
 OAI21xp33_ASAP7_75t_R n_11355 (.A1(n_11250_o_0),
    .A2(n_11353_o_0),
    .B(n_11354_o_0),
    .Y(n_11355_o_0));
 OAI31xp33_ASAP7_75t_R n_11356 (.A1(n_11223_o_0),
    .A2(n_11190_o_0),
    .A3(n_11351_o_0),
    .B(n_11355_o_0),
    .Y(n_11356_o_0));
 INVx1_ASAP7_75t_R n_11357 (.A(n_11356_o_0),
    .Y(n_11357_o_0));
 OAI211xp5_ASAP7_75t_R n_11358 (.A1(n_11189_o_0),
    .A2(n_11161_o_0),
    .B(n_11343_o_0),
    .C(n_11223_o_0),
    .Y(n_11358_o_0));
 AOI21xp33_ASAP7_75t_R n_11359 (.A1(n_11280_o_0),
    .A2(n_11345_o_0),
    .B(n_11115_o_0),
    .Y(n_11359_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1136 (.A1(n_907_o_0),
    .A2(n_887_o_0),
    .B(n_877_o_0),
    .C(n_893_o_0),
    .Y(n_1136_o_0));
 AOI21xp33_ASAP7_75t_R n_11360 (.A1(n_11276_o_0),
    .A2(n_11359_o_0),
    .B(n_11296_o_0),
    .Y(n_11360_o_0));
 AOI21xp33_ASAP7_75t_R n_11361 (.A1(n_11358_o_0),
    .A2(n_11360_o_0),
    .B(n_11192_o_0),
    .Y(n_11361_o_0));
 OAI21xp33_ASAP7_75t_R n_11362 (.A1(n_11106_o_0),
    .A2(n_11357_o_0),
    .B(n_11361_o_0),
    .Y(n_11362_o_0));
 OAI211xp5_ASAP7_75t_R n_11363 (.A1(n_11350_o_0),
    .A2(n_11224_o_0),
    .B(n_11362_o_0),
    .C(n_11220_o_0),
    .Y(n_11363_o_0));
 OAI31xp33_ASAP7_75t_R n_11364 (.A1(n_11220_o_0),
    .A2(n_11313_o_0),
    .A3(n_11333_o_0),
    .B(n_11363_o_0),
    .Y(n_11364_o_0));
 NOR2xp33_ASAP7_75t_R n_11365 (.A(n_11187_o_0),
    .B(n_11161_o_0),
    .Y(n_11365_o_0));
 AOI211xp5_ASAP7_75t_R n_11366 (.A1(n_11209_o_0),
    .A2(n_11318_o_0),
    .B(n_11365_o_0),
    .C(n_11192_o_0),
    .Y(n_11366_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11367 (.A1(net65),
    .A2(net37),
    .B(n_11250_o_0),
    .C(n_11190_o_0),
    .Y(n_11367_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11368 (.A1(n_11277_o_0),
    .A2(net65),
    .B(n_11161_o_0),
    .C(n_11177_o_1),
    .Y(n_11368_o_0));
 OAI21xp33_ASAP7_75t_R n_11369 (.A1(n_11367_o_0),
    .A2(n_11368_o_0),
    .B(n_11115_o_0),
    .Y(n_11369_o_0));
 OA21x2_ASAP7_75t_R n_1137 (.A1(n_883_o_0),
    .A2(n_1060_o_0),
    .B(n_1120_o_0),
    .Y(n_1137_o_0));
 NAND3xp33_ASAP7_75t_R n_11370 (.A(n_11136_o_0),
    .B(n_11152_o_0),
    .C(net37),
    .Y(n_11370_o_0));
 OAI211xp5_ASAP7_75t_R n_11371 (.A1(n_11186_o_0),
    .A2(net65),
    .B(n_11370_o_0),
    .C(n_11160_o_0),
    .Y(n_11371_o_0));
 OAI31xp33_ASAP7_75t_R n_11372 (.A1(n_11190_o_0),
    .A2(n_11305_o_0),
    .A3(n_11352_o_0),
    .B(n_11371_o_0),
    .Y(n_11372_o_0));
 AOI21xp33_ASAP7_75t_R n_11373 (.A1(net65),
    .A2(net37),
    .B(n_11250_o_0),
    .Y(n_11373_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11374 (.A1(n_11200_o_0),
    .A2(n_11373_o_0),
    .B(n_11265_o_0),
    .C(n_11202_o_0),
    .D(n_11223_o_0),
    .Y(n_11374_o_0));
 OAI21xp33_ASAP7_75t_R n_11375 (.A1(n_11224_o_0),
    .A2(n_11372_o_0),
    .B(n_11374_o_0),
    .Y(n_11375_o_0));
 OA21x2_ASAP7_75t_R n_11376 (.A1(n_11366_o_0),
    .A2(n_11369_o_0),
    .B(n_11375_o_0),
    .Y(n_11376_o_0));
 NAND2xp33_ASAP7_75t_R n_11377 (.A(n_11186_o_0),
    .B(n_11162_o_0),
    .Y(n_11377_o_0));
 NOR2xp33_ASAP7_75t_R n_11378 (.A(n_11251_o_0),
    .B(n_11260_o_0),
    .Y(n_11378_o_0));
 AOI31xp33_ASAP7_75t_R n_11379 (.A1(n_11165_o_0),
    .A2(n_11243_o_0),
    .A3(n_11377_o_0),
    .B(n_11378_o_0),
    .Y(n_11379_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1138 (.A1(net16),
    .A2(n_1136_o_0),
    .B(n_1137_o_0),
    .C(n_903_o_0),
    .Y(n_1138_o_0));
 AOI31xp33_ASAP7_75t_R n_11380 (.A1(n_11165_o_0),
    .A2(n_11323_o_0),
    .A3(n_11324_o_0),
    .B(n_11192_o_0),
    .Y(n_11380_o_0));
 OAI21xp33_ASAP7_75t_R n_11381 (.A1(n_11200_o_0),
    .A2(n_11351_o_0),
    .B(n_11380_o_0),
    .Y(n_11381_o_0));
 OAI21xp33_ASAP7_75t_R n_11382 (.A1(n_11202_o_0),
    .A2(n_11379_o_0),
    .B(n_11381_o_0),
    .Y(n_11382_o_0));
 INVx1_ASAP7_75t_R n_11383 (.A(n_11259_o_0),
    .Y(n_11383_o_0));
 NOR2xp33_ASAP7_75t_R n_11384 (.A(n_11136_o_0),
    .B(n_11162_o_0),
    .Y(n_11384_o_0));
 AOI31xp33_ASAP7_75t_R n_11385 (.A1(n_11160_o_0),
    .A2(n_11243_o_0),
    .A3(n_11324_o_0),
    .B(n_11224_o_0),
    .Y(n_11385_o_0));
 OAI21xp33_ASAP7_75t_R n_11386 (.A1(n_11383_o_0),
    .A2(n_11384_o_0),
    .B(n_11385_o_0),
    .Y(n_11386_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11387 (.A1(n_11207_o_0),
    .A2(n_11196_o_0),
    .B(n_11162_o_0),
    .C(n_11200_o_0),
    .Y(n_11387_o_0));
 AOI31xp33_ASAP7_75t_R n_11388 (.A1(n_11162_o_0),
    .A2(n_11190_o_0),
    .A3(net35),
    .B(n_11177_o_1),
    .Y(n_11388_o_0));
 OAI21xp33_ASAP7_75t_R n_11389 (.A1(n_11229_o_0),
    .A2(n_11387_o_0),
    .B(n_11388_o_0),
    .Y(n_11389_o_0));
 OAI211xp5_ASAP7_75t_R n_1139 (.A1(n_1133_o_0),
    .A2(n_1135_o_0),
    .B(n_930_o_0),
    .C(n_1138_o_0),
    .Y(n_1139_o_0));
 AOI31xp33_ASAP7_75t_R n_11390 (.A1(n_11223_o_0),
    .A2(n_11386_o_0),
    .A3(n_11389_o_0),
    .B(n_11220_o_0),
    .Y(n_11390_o_0));
 OAI21xp33_ASAP7_75t_R n_11391 (.A1(n_11115_o_0),
    .A2(n_11382_o_0),
    .B(n_11390_o_0),
    .Y(n_11391_o_0));
 OAI21xp33_ASAP7_75t_R n_11392 (.A1(n_11221_o_0),
    .A2(n_11376_o_0),
    .B(n_11391_o_0),
    .Y(n_11392_o_0));
 INVx1_ASAP7_75t_R n_11393 (.A(n_11296_o_0),
    .Y(n_11393_o_0));
 AOI31xp33_ASAP7_75t_R n_11394 (.A1(net35),
    .A2(net65),
    .A3(n_11190_o_0),
    .B(n_11202_o_0),
    .Y(n_11394_o_0));
 NAND2xp33_ASAP7_75t_R n_11395 (.A(n_11324_o_0),
    .B(n_11346_o_0),
    .Y(n_11395_o_0));
 AOI21xp33_ASAP7_75t_R n_11396 (.A1(n_11394_o_0),
    .A2(n_11395_o_0),
    .B(n_11115_o_0),
    .Y(n_11396_o_0));
 AOI21xp33_ASAP7_75t_R n_11397 (.A1(n_11245_o_0),
    .A2(n_11200_o_0),
    .B(n_11289_o_0),
    .Y(n_11397_o_0));
 NAND2xp33_ASAP7_75t_R n_11398 (.A(n_11202_o_0),
    .B(n_11397_o_0),
    .Y(n_11398_o_0));
 INVx1_ASAP7_75t_R n_11399 (.A(n_11201_o_0),
    .Y(n_11399_o_0));
 OAI21xp33_ASAP7_75t_R n_1140 (.A1(n_847_o_0),
    .A2(net32),
    .B(n_1121_o_0),
    .Y(n_1140_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11400 (.A1(n_11264_o_0),
    .A2(net65),
    .B(n_11276_o_0),
    .C(n_11202_o_0),
    .Y(n_11400_o_0));
 AOI21xp33_ASAP7_75t_R n_11401 (.A1(n_11160_o_0),
    .A2(n_11399_o_0),
    .B(n_11400_o_0),
    .Y(n_11401_o_0));
 OAI21xp33_ASAP7_75t_R n_11402 (.A1(net58),
    .A2(net65),
    .B(n_11200_o_0),
    .Y(n_11402_o_0));
 INVx1_ASAP7_75t_R n_11403 (.A(n_11179_o_0),
    .Y(n_11403_o_0));
 OAI21xp33_ASAP7_75t_R n_11404 (.A1(n_11402_o_0),
    .A2(n_11403_o_0),
    .B(n_11192_o_0),
    .Y(n_11404_o_0));
 AOI21xp33_ASAP7_75t_R n_11405 (.A1(n_11354_o_0),
    .A2(n_11268_o_0),
    .B(n_11404_o_0),
    .Y(n_11405_o_0));
 OAI31xp33_ASAP7_75t_R n_11406 (.A1(n_11212_o_0),
    .A2(n_11401_o_0),
    .A3(n_11405_o_0),
    .B(n_11221_o_0),
    .Y(n_11406_o_0));
 OAI21xp33_ASAP7_75t_R n_11407 (.A1(n_11159_o_0),
    .A2(n_11199_o_0),
    .B(n_11162_o_0),
    .Y(n_11407_o_0));
 OAI21xp33_ASAP7_75t_R n_11408 (.A1(n_11159_o_0),
    .A2(n_11199_o_0),
    .B(n_11152_o_0),
    .Y(n_11408_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11409 (.A1(n_11196_o_0),
    .A2(n_11207_o_0),
    .B(n_11407_o_0),
    .C(n_11408_o_0),
    .D(n_11384_o_0),
    .Y(n_11409_o_0));
 OAI31xp33_ASAP7_75t_R n_1141 (.A1(n_878_o_0),
    .A2(n_1050_o_0),
    .A3(n_945_o_0),
    .B(n_1140_o_0),
    .Y(n_1141_o_0));
 AOI31xp33_ASAP7_75t_R n_11410 (.A1(n_11165_o_0),
    .A2(n_11195_o_0),
    .A3(n_11353_o_0),
    .B(n_11409_o_0),
    .Y(n_11410_o_0));
 NOR2xp33_ASAP7_75t_R n_11411 (.A(n_11152_o_0),
    .B(n_11277_o_0),
    .Y(n_11411_o_0));
 NAND2xp33_ASAP7_75t_R n_11412 (.A(n_11200_o_0),
    .B(n_11179_o_0),
    .Y(n_11412_o_0));
 OAI211xp5_ASAP7_75t_R n_11413 (.A1(n_11411_o_0),
    .A2(n_11412_o_0),
    .B(n_11290_o_0),
    .C(n_11224_o_0),
    .Y(n_11413_o_0));
 OAI21xp33_ASAP7_75t_R n_11414 (.A1(n_11202_o_0),
    .A2(n_11410_o_0),
    .B(n_11413_o_0),
    .Y(n_11414_o_0));
 OAI21xp33_ASAP7_75t_R n_11415 (.A1(net68),
    .A2(n_11250_o_0),
    .B(n_11152_o_0),
    .Y(n_11415_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11416 (.A1(n_11152_o_0),
    .A2(n_11282_o_0),
    .B(n_11415_o_0),
    .C(n_11190_o_0),
    .Y(n_11416_o_0));
 AOI31xp33_ASAP7_75t_R n_11417 (.A1(n_11160_o_0),
    .A2(n_11243_o_0),
    .A3(n_11324_o_0),
    .B(n_11416_o_0),
    .Y(n_11417_o_0));
 OAI21xp33_ASAP7_75t_R n_11418 (.A1(n_11139_o_0),
    .A2(n_11250_o_0),
    .B(n_11152_o_0),
    .Y(n_11418_o_0));
 INVx1_ASAP7_75t_R n_11419 (.A(n_11418_o_0),
    .Y(n_11419_o_0));
 NAND2xp33_ASAP7_75t_R n_1142 (.A(n_878_o_0),
    .B(n_982_o_0),
    .Y(n_1142_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11420 (.A1(n_11328_o_0),
    .A2(n_11419_o_0),
    .B(n_11395_o_0),
    .C(n_11224_o_0),
    .Y(n_11420_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11421 (.A1(n_11202_o_0),
    .A2(n_11417_o_0),
    .B(n_11420_o_0),
    .C(n_11266_o_0),
    .D(n_11221_o_0),
    .Y(n_11421_o_0));
 OAI21xp33_ASAP7_75t_R n_11422 (.A1(n_11212_o_0),
    .A2(n_11414_o_0),
    .B(n_11421_o_0),
    .Y(n_11422_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11423 (.A1(n_11396_o_0),
    .A2(n_11398_o_0),
    .B(n_11406_o_0),
    .C(n_11422_o_0),
    .Y(n_11423_o_0));
 OAI22xp33_ASAP7_75t_R n_11424 (.A1(n_11392_o_0),
    .A2(n_11105_o_0),
    .B1(n_11393_o_0),
    .B2(n_11423_o_0),
    .Y(n_11424_o_0));
 NAND2xp33_ASAP7_75t_R n_11425 (.A(net65),
    .B(n_11264_o_0),
    .Y(n_11425_o_0));
 AOI31xp33_ASAP7_75t_R n_11426 (.A1(n_11165_o_0),
    .A2(n_11292_o_0),
    .A3(n_11425_o_0),
    .B(n_11409_o_0),
    .Y(n_11426_o_0));
 OAI21xp33_ASAP7_75t_R n_11427 (.A1(net49),
    .A2(n_11426_o_0),
    .B(n_11296_o_0),
    .Y(n_11427_o_0));
 AO21x1_ASAP7_75t_R n_11428 (.A1(n_11377_o_0),
    .A2(n_11306_o_0),
    .B(n_11224_o_0),
    .Y(n_11428_o_0));
 AOI21xp33_ASAP7_75t_R n_11429 (.A1(n_11240_o_0),
    .A2(n_11209_o_0),
    .B(n_11428_o_0),
    .Y(n_11429_o_0));
 OAI31xp33_ASAP7_75t_R n_1143 (.A1(n_878_o_0),
    .A2(n_934_o_0),
    .A3(n_1006_o_0),
    .B(n_1142_o_0),
    .Y(n_1143_o_0));
 AOI21xp33_ASAP7_75t_R n_11430 (.A1(n_11152_o_0),
    .A2(n_11197_o_0),
    .B(n_11200_o_0),
    .Y(n_11430_o_0));
 OA21x2_ASAP7_75t_R n_11431 (.A1(net65),
    .A2(n_11186_o_0),
    .B(n_11346_o_0),
    .Y(n_11431_o_0));
 AOI21xp33_ASAP7_75t_R n_11432 (.A1(n_11430_o_0),
    .A2(n_11345_o_0),
    .B(n_11431_o_0),
    .Y(n_11432_o_0));
 OAI21xp33_ASAP7_75t_R n_11433 (.A1(n_11162_o_0),
    .A2(n_11187_o_0),
    .B(n_11185_o_0),
    .Y(n_11433_o_0));
 AOI21xp33_ASAP7_75t_R n_11434 (.A1(n_11433_o_0),
    .A2(n_11178_o_0),
    .B(n_11105_o_0),
    .Y(n_11434_o_0));
 OAI21xp33_ASAP7_75t_R n_11435 (.A1(net49),
    .A2(n_11432_o_0),
    .B(n_11434_o_0),
    .Y(n_11435_o_0));
 OAI211xp5_ASAP7_75t_R n_11436 (.A1(n_11427_o_0),
    .A2(n_11429_o_0),
    .B(n_11115_o_0),
    .C(n_11435_o_0),
    .Y(n_11436_o_0));
 AOI21xp33_ASAP7_75t_R n_11437 (.A1(n_11393_o_0),
    .A2(n_11346_o_0),
    .B(n_11192_o_0),
    .Y(n_11437_o_0));
 OAI21xp33_ASAP7_75t_R n_11438 (.A1(n_11172_o_0),
    .A2(n_11161_o_0),
    .B(n_11437_o_0),
    .Y(n_11438_o_0));
 NOR3xp33_ASAP7_75t_R n_11439 (.A(n_11276_o_0),
    .B(n_11384_o_0),
    .C(n_11106_o_0),
    .Y(n_11439_o_0));
 OA21x2_ASAP7_75t_R n_1144 (.A1(n_1143_o_0),
    .A2(net42),
    .B(n_904_o_0),
    .Y(n_1144_o_0));
 NAND3xp33_ASAP7_75t_R n_11440 (.A(n_11197_o_0),
    .B(n_11165_o_0),
    .C(net65),
    .Y(n_11440_o_0));
 OAI21xp33_ASAP7_75t_R n_11441 (.A1(n_11161_o_0),
    .A2(n_11341_o_0),
    .B(n_11440_o_0),
    .Y(n_11441_o_0));
 NAND2xp33_ASAP7_75t_R n_11442 (.A(n_11152_o_0),
    .B(n_11186_o_0),
    .Y(n_11442_o_0));
 OAI211xp5_ASAP7_75t_R n_11443 (.A1(n_11197_o_0),
    .A2(net65),
    .B(n_11160_o_0),
    .C(n_11442_o_0),
    .Y(n_11443_o_0));
 OAI31xp33_ASAP7_75t_R n_11444 (.A1(n_11190_o_0),
    .A2(n_11278_o_0),
    .A3(n_11314_o_0),
    .B(n_11443_o_0),
    .Y(n_11444_o_0));
 AOI21xp33_ASAP7_75t_R n_11445 (.A1(n_11393_o_0),
    .A2(n_11444_o_0),
    .B(n_11224_o_0),
    .Y(n_11445_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11446 (.A1(n_11106_o_0),
    .A2(n_11441_o_0),
    .B(n_11445_o_0),
    .C(n_11223_o_0),
    .Y(n_11446_o_0));
 OAI21xp33_ASAP7_75t_R n_11447 (.A1(n_11438_o_0),
    .A2(n_11439_o_0),
    .B(n_11446_o_0),
    .Y(n_11447_o_0));
 NAND2xp33_ASAP7_75t_R n_11448 (.A(n_11162_o_0),
    .B(n_11187_o_0),
    .Y(n_11448_o_0));
 AOI21xp33_ASAP7_75t_R n_11449 (.A1(n_11165_o_0),
    .A2(n_11448_o_0),
    .B(n_11365_o_0),
    .Y(n_11449_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1145 (.A1(net16),
    .A2(n_1141_o_0),
    .B(n_903_o_0),
    .C(n_1144_o_0),
    .Y(n_1145_o_0));
 NAND2xp33_ASAP7_75t_R n_11450 (.A(n_11139_o_0),
    .B(n_11152_o_0),
    .Y(n_11450_o_0));
 AOI21xp33_ASAP7_75t_R n_11451 (.A1(n_11450_o_0),
    .A2(n_11185_o_0),
    .B(n_11223_o_0),
    .Y(n_11451_o_0));
 OAI21xp33_ASAP7_75t_R n_11452 (.A1(n_11402_o_0),
    .A2(n_11419_o_0),
    .B(n_11451_o_0),
    .Y(n_11452_o_0));
 OAI21xp33_ASAP7_75t_R n_11453 (.A1(n_11266_o_0),
    .A2(n_11449_o_0),
    .B(n_11452_o_0),
    .Y(n_11453_o_0));
 NOR2xp33_ASAP7_75t_R n_11454 (.A(n_11152_o_0),
    .B(n_11165_o_0),
    .Y(n_11454_o_0));
 NAND2xp33_ASAP7_75t_R n_11455 (.A(n_11197_o_0),
    .B(n_11454_o_0),
    .Y(n_11455_o_0));
 NAND2xp33_ASAP7_75t_R n_11456 (.A(net65),
    .B(n_11165_o_0),
    .Y(n_11456_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11457 (.A1(n_11196_o_0),
    .A2(n_11207_o_0),
    .B(n_11456_o_0),
    .C(n_11266_o_0),
    .Y(n_11457_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11458 (.A1(net35),
    .A2(n_11162_o_0),
    .B(n_11354_o_0),
    .C(n_11324_o_0),
    .D(n_11457_o_0),
    .Y(n_11458_o_0));
 AOI211xp5_ASAP7_75t_R n_11459 (.A1(n_11115_o_0),
    .A2(n_11455_o_0),
    .B(n_11458_o_0),
    .C(n_11296_o_0),
    .Y(n_11459_o_0));
 NOR2xp33_ASAP7_75t_R n_1146 (.A(n_881_o_0),
    .B(n_918_o_0),
    .Y(n_1146_o_0));
 INVx1_ASAP7_75t_R n_11460 (.A(n_11324_o_0),
    .Y(n_11460_o_0));
 OAI211xp5_ASAP7_75t_R n_11461 (.A1(n_11230_o_0),
    .A2(n_11460_o_0),
    .B(n_11440_o_0),
    .C(n_11266_o_0),
    .Y(n_11461_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11462 (.A1(n_11188_o_0),
    .A2(n_11231_o_0),
    .B(n_11192_o_0),
    .C(n_11393_o_0),
    .Y(n_11462_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11463 (.A1(n_11197_o_0),
    .A2(n_11454_o_0),
    .B(n_11266_o_0),
    .C(n_11461_o_0),
    .D(n_11462_o_0),
    .Y(n_11463_o_0));
 AOI211xp5_ASAP7_75t_R n_11464 (.A1(n_11453_o_0),
    .A2(n_11224_o_0),
    .B(n_11459_o_0),
    .C(n_11463_o_0),
    .Y(n_11464_o_0));
 INVx1_ASAP7_75t_R n_11465 (.A(n_11442_o_0),
    .Y(n_11465_o_0));
 NOR2xp33_ASAP7_75t_R n_11466 (.A(n_11139_o_0),
    .B(n_11152_o_0),
    .Y(n_11466_o_0));
 OAI31xp33_ASAP7_75t_R n_11467 (.A1(n_11190_o_0),
    .A2(n_11465_o_0),
    .A3(n_11466_o_0),
    .B(n_11355_o_0),
    .Y(n_11467_o_0));
 AOI21xp33_ASAP7_75t_R n_11468 (.A1(n_11224_o_0),
    .A2(n_11467_o_0),
    .B(n_11115_o_0),
    .Y(n_11468_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11469 (.A1(n_11188_o_0),
    .A2(n_11162_o_0),
    .B(n_11329_o_0),
    .C(n_11200_o_0),
    .Y(n_11469_o_0));
 NOR4xp25_ASAP7_75t_R n_1147 (.A(n_1146_o_0),
    .B(n_989_o_0),
    .C(n_904_o_0),
    .D(n_878_o_0),
    .Y(n_1147_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11470 (.A1(n_11260_o_0),
    .A2(n_11137_o_0),
    .B(n_11469_o_0),
    .C(n_11192_o_0),
    .Y(n_11470_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11471 (.A1(n_11186_o_0),
    .A2(n_11152_o_0),
    .B(n_11327_o_0),
    .C(n_11160_o_0),
    .Y(n_11471_o_0));
 AOI21xp33_ASAP7_75t_R n_11472 (.A1(n_11418_o_0),
    .A2(n_11185_o_0),
    .B(n_11471_o_0),
    .Y(n_11472_o_0));
 INVx1_ASAP7_75t_R n_11473 (.A(n_11114_o_0),
    .Y(n_11473_o_0));
 NOR2xp33_ASAP7_75t_R n_11474 (.A(n_11113_o_0),
    .B(n_11112_o_0),
    .Y(n_11474_o_0));
 OAI22xp33_ASAP7_75t_R n_11475 (.A1(n_11472_o_0),
    .A2(n_11224_o_0),
    .B1(n_11473_o_0),
    .B2(n_11474_o_0),
    .Y(n_11475_o_0));
 OAI21xp33_ASAP7_75t_R n_11476 (.A1(n_11470_o_0),
    .A2(n_11475_o_0),
    .B(n_11106_o_0),
    .Y(n_11476_o_0));
 AOI21xp33_ASAP7_75t_R n_11477 (.A1(n_11368_o_0),
    .A2(n_11468_o_0),
    .B(n_11476_o_0),
    .Y(n_11477_o_0));
 OAI21xp33_ASAP7_75t_R n_11478 (.A1(n_11464_o_0),
    .A2(n_11477_o_0),
    .B(n_11220_o_0),
    .Y(n_11478_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11479 (.A1(n_11436_o_0),
    .A2(n_11447_o_0),
    .B(n_11220_o_0),
    .C(n_11478_o_0),
    .Y(n_11479_o_0));
 NAND3xp33_ASAP7_75t_R n_1148 (.A(n_889_o_0),
    .B(n_881_o_0),
    .C(n_877_o_0),
    .Y(n_1148_o_0));
 AO21x1_ASAP7_75t_R n_11480 (.A1(n_11197_o_0),
    .A2(net65),
    .B(n_11334_o_0),
    .Y(n_11480_o_0));
 AOI21xp33_ASAP7_75t_R n_11481 (.A1(n_11206_o_0),
    .A2(n_11240_o_0),
    .B(n_11160_o_0),
    .Y(n_11481_o_0));
 NOR3xp33_ASAP7_75t_R n_11482 (.A(n_11236_o_0),
    .B(n_11481_o_0),
    .C(n_11223_o_0),
    .Y(n_11482_o_0));
 AOI31xp33_ASAP7_75t_R n_11483 (.A1(n_11228_o_0),
    .A2(n_11115_o_0),
    .A3(n_11480_o_0),
    .B(n_11482_o_0),
    .Y(n_11483_o_0));
 NOR2xp33_ASAP7_75t_R n_11484 (.A(n_11328_o_0),
    .B(n_11419_o_0),
    .Y(n_11484_o_0));
 AOI211xp5_ASAP7_75t_R n_11485 (.A1(net65),
    .A2(n_11250_o_0),
    .B(n_11229_o_0),
    .C(n_11160_o_0),
    .Y(n_11485_o_0));
 NAND4xp25_ASAP7_75t_R n_11486 (.A(n_11207_o_0),
    .B(n_11196_o_0),
    .C(net65),
    .D(n_11200_o_0),
    .Y(n_11486_o_0));
 NAND4xp25_ASAP7_75t_R n_11487 (.A(n_11486_o_0),
    .B(n_11448_o_0),
    .C(n_11267_o_0),
    .D(n_11115_o_0),
    .Y(n_11487_o_0));
 OAI31xp33_ASAP7_75t_R n_11488 (.A1(n_11223_o_0),
    .A2(n_11484_o_0),
    .A3(n_11485_o_0),
    .B(n_11487_o_0),
    .Y(n_11488_o_0));
 OAI21xp33_ASAP7_75t_R n_11489 (.A1(n_11224_o_0),
    .A2(n_11488_o_0),
    .B(n_11105_o_0),
    .Y(n_11489_o_0));
 OAI32xp33_ASAP7_75t_R n_1149 (.A1(n_881_o_0),
    .A2(n_1061_o_0),
    .A3(n_1044_o_0),
    .B1(n_1148_o_0),
    .B2(n_903_o_0),
    .Y(n_1149_o_0));
 AOI21xp33_ASAP7_75t_R n_11490 (.A1(n_11202_o_0),
    .A2(n_11483_o_0),
    .B(n_11489_o_0),
    .Y(n_11490_o_0));
 INVx1_ASAP7_75t_R n_11491 (.A(n_11342_o_0),
    .Y(n_11491_o_0));
 NAND3xp33_ASAP7_75t_R n_11492 (.A(n_11323_o_0),
    .B(n_11324_o_0),
    .C(n_11165_o_0),
    .Y(n_11492_o_0));
 OAI21xp33_ASAP7_75t_R n_11493 (.A1(n_11274_o_0),
    .A2(n_11189_o_0),
    .B(n_11223_o_0),
    .Y(n_11493_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11494 (.A1(n_11206_o_0),
    .A2(n_11259_o_0),
    .B(n_11493_o_0),
    .C(n_11224_o_0),
    .Y(n_11494_o_0));
 NOR3xp33_ASAP7_75t_R n_11495 (.A(n_11189_o_0),
    .B(n_11314_o_0),
    .C(n_11190_o_0),
    .Y(n_11495_o_0));
 NAND2xp33_ASAP7_75t_R n_11496 (.A(n_11152_o_0),
    .B(n_11250_o_0),
    .Y(n_11496_o_0));
 AOI21xp33_ASAP7_75t_R n_11497 (.A1(n_11282_o_0),
    .A2(n_11496_o_0),
    .B(n_11165_o_0),
    .Y(n_11497_o_0));
 AOI21xp33_ASAP7_75t_R n_11498 (.A1(n_11165_o_0),
    .A2(n_11442_o_0),
    .B(n_11212_o_0),
    .Y(n_11498_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11499 (.A1(n_11188_o_0),
    .A2(net65),
    .B(n_11498_o_0),
    .C(n_11202_o_0),
    .Y(n_11499_o_0));
 INVx1_ASAP7_75t_R n_1150 (.A(n_1001_o_0),
    .Y(n_1150_o_0));
 OAI31xp33_ASAP7_75t_R n_11500 (.A1(n_11223_o_0),
    .A2(n_11495_o_0),
    .A3(n_11497_o_0),
    .B(n_11499_o_0),
    .Y(n_11500_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11501 (.A1(n_11491_o_0),
    .A2(n_11492_o_0),
    .B(n_11494_o_0),
    .C(n_11500_o_0),
    .Y(n_11501_o_0));
 NOR2xp33_ASAP7_75t_R n_11502 (.A(n_11105_o_0),
    .B(n_11501_o_0),
    .Y(n_11502_o_0));
 NAND2xp33_ASAP7_75t_R n_11503 (.A(n_11152_o_0),
    .B(n_11250_o_0),
    .Y(n_11503_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11504 (.A1(n_11201_o_0),
    .A2(n_11503_o_0),
    .B(n_11200_o_0),
    .C(n_11343_o_0),
    .Y(n_11504_o_0));
 INVx1_ASAP7_75t_R n_11505 (.A(n_11504_o_0),
    .Y(n_11505_o_0));
 OAI21xp33_ASAP7_75t_R n_11506 (.A1(n_11161_o_0),
    .A2(n_11278_o_0),
    .B(n_11202_o_0),
    .Y(n_11506_o_0));
 AOI21xp33_ASAP7_75t_R n_11507 (.A1(net65),
    .A2(n_11165_o_0),
    .B(n_11506_o_0),
    .Y(n_11507_o_0));
 AOI211xp5_ASAP7_75t_R n_11508 (.A1(net49),
    .A2(n_11505_o_0),
    .B(n_11507_o_0),
    .C(n_11223_o_0),
    .Y(n_11508_o_0));
 INVx1_ASAP7_75t_R n_11509 (.A(n_11412_o_0),
    .Y(n_11509_o_0));
 NOR4xp25_ASAP7_75t_R n_1151 (.A(n_1147_o_0),
    .B(n_1149_o_0),
    .C(net14),
    .D(n_1150_o_0),
    .Y(n_1151_o_0));
 AOI21xp33_ASAP7_75t_R n_11510 (.A1(net65),
    .A2(n_11188_o_0),
    .B(n_11165_o_0),
    .Y(n_11510_o_0));
 INVx1_ASAP7_75t_R n_11511 (.A(n_11197_o_0),
    .Y(n_11511_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11512 (.A1(net65),
    .A2(n_11511_o_0),
    .B(n_11328_o_0),
    .C(n_11270_o_0),
    .Y(n_11512_o_0));
 OAI31xp33_ASAP7_75t_R n_11513 (.A1(n_11202_o_0),
    .A2(n_11509_o_0),
    .A3(n_11510_o_0),
    .B(n_11512_o_0),
    .Y(n_11513_o_0));
 OAI21xp33_ASAP7_75t_R n_11514 (.A1(n_11212_o_0),
    .A2(n_11513_o_0),
    .B(n_11393_o_0),
    .Y(n_11514_o_0));
 NOR2xp33_ASAP7_75t_R n_11515 (.A(n_11172_o_0),
    .B(n_11166_o_0),
    .Y(n_11515_o_0));
 OAI211xp5_ASAP7_75t_R n_11516 (.A1(n_11190_o_0),
    .A2(net65),
    .B(n_11250_o_0),
    .C(net37),
    .Y(n_11516_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11517 (.A1(n_11162_o_0),
    .A2(net58),
    .B(n_11190_o_0),
    .C(n_11186_o_0),
    .Y(n_11517_o_0));
 AOI211xp5_ASAP7_75t_R n_11518 (.A1(n_11516_o_0),
    .A2(n_11517_o_0),
    .B(n_11497_o_0),
    .C(n_11202_o_0),
    .Y(n_11518_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11519 (.A1(n_11515_o_0),
    .A2(n_11253_o_0),
    .B(n_11224_o_0),
    .C(n_11518_o_0),
    .Y(n_11519_o_0));
 NOR3xp33_ASAP7_75t_R n_1152 (.A(n_1006_o_0),
    .B(n_877_o_0),
    .C(n_907_o_0),
    .Y(n_1152_o_0));
 OAI211xp5_ASAP7_75t_R n_11520 (.A1(net35),
    .A2(n_11152_o_0),
    .B(n_11442_o_0),
    .C(n_11165_o_0),
    .Y(n_11520_o_0));
 OAI21xp33_ASAP7_75t_R n_11521 (.A1(n_11172_o_0),
    .A2(n_11407_o_0),
    .B(n_11520_o_0),
    .Y(n_11521_o_0));
 NOR2xp33_ASAP7_75t_R n_11522 (.A(n_11162_o_0),
    .B(n_11160_o_0),
    .Y(n_11522_o_0));
 OAI21xp33_ASAP7_75t_R n_11523 (.A1(n_11165_o_0),
    .A2(n_11291_o_0),
    .B(n_11224_o_0),
    .Y(n_11523_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11524 (.A1(n_11511_o_0),
    .A2(n_11522_o_0),
    .B(n_11523_o_0),
    .C(n_11223_o_0),
    .Y(n_11524_o_0));
 AOI21xp33_ASAP7_75t_R n_11525 (.A1(n_11192_o_0),
    .A2(n_11521_o_0),
    .B(n_11524_o_0),
    .Y(n_11525_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11526 (.A1(n_11519_o_0),
    .A2(n_11266_o_0),
    .B(n_11525_o_0),
    .C(n_11296_o_0),
    .Y(n_11526_o_0));
 OAI211xp5_ASAP7_75t_R n_11527 (.A1(n_11508_o_0),
    .A2(n_11514_o_0),
    .B(n_11526_o_0),
    .C(n_11220_o_0),
    .Y(n_11527_o_0));
 OAI31xp33_ASAP7_75t_R n_11528 (.A1(n_11220_o_0),
    .A2(n_11490_o_0),
    .A3(n_11502_o_0),
    .B(n_11527_o_0),
    .Y(n_11528_o_0));
 OAI311xp33_ASAP7_75t_R n_11529 (.A1(n_11190_o_0),
    .A2(n_11172_o_0),
    .A3(n_11162_o_0),
    .B1(n_11177_o_1),
    .C1(n_11328_o_0),
    .Y(n_11529_o_0));
 INVx1_ASAP7_75t_R n_1153 (.A(n_1152_o_0),
    .Y(n_1153_o_0));
 OAI31xp33_ASAP7_75t_R n_11530 (.A1(net49),
    .A2(n_11471_o_0),
    .A3(n_11185_o_0),
    .B(n_11529_o_0),
    .Y(n_11530_o_0));
 INVx1_ASAP7_75t_R n_11531 (.A(n_11530_o_0),
    .Y(n_11531_o_0));
 NAND2xp33_ASAP7_75t_R n_11532 (.A(net35),
    .B(n_11162_o_0),
    .Y(n_11532_o_0));
 AOI22xp33_ASAP7_75t_R n_11533 (.A1(n_11511_o_0),
    .A2(n_11522_o_0),
    .B1(n_11532_o_0),
    .B2(n_11510_o_0),
    .Y(n_11533_o_0));
 AOI21xp33_ASAP7_75t_R n_11534 (.A1(n_11160_o_0),
    .A2(n_11370_o_0),
    .B(n_11192_o_0),
    .Y(n_11534_o_0));
 OAI21xp33_ASAP7_75t_R n_11535 (.A1(n_11251_o_0),
    .A2(n_11276_o_0),
    .B(n_11534_o_0),
    .Y(n_11535_o_0));
 OAI211xp5_ASAP7_75t_R n_11536 (.A1(n_11533_o_0),
    .A2(n_11224_o_0),
    .B(n_11535_o_0),
    .C(n_11105_o_0),
    .Y(n_11536_o_0));
 OAI21xp33_ASAP7_75t_R n_11537 (.A1(n_11296_o_0),
    .A2(n_11531_o_0),
    .B(n_11536_o_0),
    .Y(n_11537_o_0));
 NAND3xp33_ASAP7_75t_R n_11538 (.A(n_11309_o_0),
    .B(n_11327_o_0),
    .C(n_11160_o_0),
    .Y(n_11538_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11539 (.A1(n_11258_o_0),
    .A2(n_11345_o_0),
    .B(n_11160_o_0),
    .C(n_11538_o_0),
    .Y(n_11539_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1154 (.A1(n_1153_o_0),
    .A2(n_1062_o_0),
    .B(net16),
    .C(n_1079_o_0),
    .Y(n_1154_o_0));
 AOI211xp5_ASAP7_75t_R n_11540 (.A1(net35),
    .A2(n_11200_o_0),
    .B(n_11497_o_0),
    .C(n_11177_o_1),
    .Y(n_11540_o_0));
 AOI21xp33_ASAP7_75t_R n_11541 (.A1(n_11192_o_0),
    .A2(n_11539_o_0),
    .B(n_11540_o_0),
    .Y(n_11541_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11542 (.A1(n_11136_o_0),
    .A2(net37),
    .B(n_11162_o_0),
    .C(n_11200_o_0),
    .Y(n_11542_o_0));
 AOI21xp33_ASAP7_75t_R n_11543 (.A1(n_11162_o_0),
    .A2(n_11264_o_0),
    .B(n_11542_o_0),
    .Y(n_11543_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11544 (.A1(n_11250_o_0),
    .A2(net37),
    .B(n_11162_o_0),
    .C(n_11190_o_0),
    .Y(n_11544_o_0));
 OAI321xp33_ASAP7_75t_R n_11545 (.A1(net37),
    .A2(n_11235_o_0),
    .A3(n_11160_o_0),
    .B1(n_11229_o_0),
    .B2(n_11544_o_0),
    .C(n_11192_o_0),
    .Y(n_11545_o_0));
 OAI31xp33_ASAP7_75t_R n_11546 (.A1(net49),
    .A2(n_11286_o_0),
    .A3(n_11543_o_0),
    .B(n_11545_o_0),
    .Y(n_11546_o_0));
 AOI21xp33_ASAP7_75t_R n_11547 (.A1(n_11393_o_0),
    .A2(n_11546_o_0),
    .B(n_11212_o_0),
    .Y(n_11547_o_0));
 OAI21xp33_ASAP7_75t_R n_11548 (.A1(n_11106_o_0),
    .A2(n_11541_o_0),
    .B(n_11547_o_0),
    .Y(n_11548_o_0));
 OAI21xp33_ASAP7_75t_R n_11549 (.A1(n_11223_o_0),
    .A2(n_11537_o_0),
    .B(n_11548_o_0),
    .Y(n_11549_o_0));
 NOR2xp33_ASAP7_75t_R n_1155 (.A(n_933_o_0),
    .B(n_881_o_0),
    .Y(n_1155_o_0));
 INVx1_ASAP7_75t_R n_11550 (.A(n_11327_o_0),
    .Y(n_11550_o_0));
 INVx1_ASAP7_75t_R n_11551 (.A(n_11345_o_0),
    .Y(n_11551_o_0));
 AO21x1_ASAP7_75t_R n_11552 (.A1(n_11264_o_0),
    .A2(net65),
    .B(n_11274_o_0),
    .Y(n_11552_o_0));
 OAI31xp33_ASAP7_75t_R n_11553 (.A1(n_11190_o_0),
    .A2(n_11550_o_0),
    .A3(n_11551_o_0),
    .B(n_11552_o_0),
    .Y(n_11553_o_0));
 INVx1_ASAP7_75t_R n_11554 (.A(n_11161_o_0),
    .Y(n_11554_o_0));
 AOI21xp33_ASAP7_75t_R n_11555 (.A1(n_11323_o_0),
    .A2(n_11554_o_0),
    .B(n_11212_o_0),
    .Y(n_11555_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11556 (.A1(net58),
    .A2(n_11190_o_0),
    .B(n_11555_o_0),
    .C(n_11177_o_1),
    .Y(n_11556_o_0));
 OAI21xp33_ASAP7_75t_R n_11557 (.A1(n_11115_o_0),
    .A2(n_11553_o_0),
    .B(n_11556_o_0),
    .Y(n_11557_o_0));
 AOI21xp33_ASAP7_75t_R n_11558 (.A1(net65),
    .A2(n_11172_o_0),
    .B(n_11276_o_0),
    .Y(n_11558_o_0));
 AOI21xp33_ASAP7_75t_R n_11559 (.A1(n_11250_o_0),
    .A2(n_11162_o_0),
    .B(n_11544_o_0),
    .Y(n_11559_o_0));
 OAI21xp33_ASAP7_75t_R n_1156 (.A1(n_982_o_0),
    .A2(n_1155_o_0),
    .B(n_878_o_0),
    .Y(n_1156_o_0));
 INVx1_ASAP7_75t_R n_11560 (.A(n_11268_o_0),
    .Y(n_11560_o_0));
 OAI321xp33_ASAP7_75t_R n_11561 (.A1(n_11419_o_0),
    .A2(n_11560_o_0),
    .A3(n_11165_o_0),
    .B1(n_11160_o_0),
    .B2(n_11442_o_0),
    .C(n_11212_o_0),
    .Y(n_11561_o_0));
 OAI311xp33_ASAP7_75t_R n_11562 (.A1(n_11266_o_0),
    .A2(n_11558_o_0),
    .A3(n_11559_o_0),
    .B1(net49),
    .C1(n_11561_o_0),
    .Y(n_11562_o_0));
 OAI21xp33_ASAP7_75t_R n_11563 (.A1(n_11152_o_0),
    .A2(n_11197_o_0),
    .B(n_11160_o_0),
    .Y(n_11563_o_0));
 OAI22xp33_ASAP7_75t_R n_11564 (.A1(n_11278_o_0),
    .A2(n_11563_o_0),
    .B1(n_11276_o_0),
    .B2(n_11257_o_0),
    .Y(n_11564_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11565 (.A1(n_11267_o_0),
    .A2(n_11542_o_0),
    .B(n_11212_o_0),
    .C(n_11192_o_0),
    .Y(n_11565_o_0));
 OAI21xp33_ASAP7_75t_R n_11566 (.A1(n_11190_o_0),
    .A2(n_11187_o_0),
    .B(n_11266_o_0),
    .Y(n_11566_o_0));
 AOI21xp33_ASAP7_75t_R n_11567 (.A1(n_11160_o_0),
    .A2(n_11345_o_0),
    .B(n_11566_o_0),
    .Y(n_11567_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11568 (.A1(net37),
    .A2(n_11162_o_0),
    .B(n_11160_o_0),
    .C(n_11115_o_0),
    .Y(n_11568_o_0));
 AOI21xp33_ASAP7_75t_R n_11569 (.A1(n_11289_o_0),
    .A2(n_11268_o_0),
    .B(n_11568_o_0),
    .Y(n_11569_o_0));
 NAND3xp33_ASAP7_75t_R n_1157 (.A(n_939_o_0),
    .B(n_882_o_0),
    .C(n_877_o_0),
    .Y(n_1157_o_0));
 OAI211xp5_ASAP7_75t_R n_11570 (.A1(n_11567_o_0),
    .A2(n_11569_o_0),
    .B(n_11224_o_0),
    .C(n_11105_o_0),
    .Y(n_11570_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11571 (.A1(n_11266_o_0),
    .A2(n_11564_o_0),
    .B(n_11565_o_0),
    .C(n_11570_o_0),
    .Y(n_11571_o_0));
 NAND2xp33_ASAP7_75t_R n_11572 (.A(net65),
    .B(n_11291_o_0),
    .Y(n_11572_o_0));
 AOI22xp33_ASAP7_75t_R n_11573 (.A1(n_11198_o_0),
    .A2(n_11258_o_0),
    .B1(n_11572_o_0),
    .B2(n_11208_o_0),
    .Y(n_11573_o_0));
 INVx1_ASAP7_75t_R n_11574 (.A(n_11565_o_0),
    .Y(n_11574_o_0));
 OAI211xp5_ASAP7_75t_R n_11575 (.A1(n_11573_o_0),
    .A2(n_11115_o_0),
    .B(n_11574_o_0),
    .C(n_11106_o_0),
    .Y(n_11575_o_0));
 AOI321xp33_ASAP7_75t_R n_11576 (.A1(n_11106_o_0),
    .A2(n_11557_o_0),
    .A3(n_11562_o_0),
    .B1(n_11571_o_0),
    .B2(n_11575_o_0),
    .C(n_11221_o_0),
    .Y(n_11576_o_0));
 AO21x1_ASAP7_75t_R n_11577 (.A1(n_11549_o_0),
    .A2(n_11221_o_0),
    .B(n_11576_o_0),
    .Y(n_11577_o_0));
 AOI21xp33_ASAP7_75t_R n_11578 (.A1(n_11370_o_0),
    .A2(n_11198_o_0),
    .B(n_11224_o_0),
    .Y(n_11578_o_0));
 OAI21xp33_ASAP7_75t_R n_11579 (.A1(n_11200_o_0),
    .A2(n_11329_o_0),
    .B(n_11578_o_0),
    .Y(n_11579_o_0));
 AOI21xp33_ASAP7_75t_R n_1158 (.A1(n_1156_o_0),
    .A2(n_1157_o_0),
    .B(n_891_o_0),
    .Y(n_1158_o_0));
 NAND2xp33_ASAP7_75t_R n_11580 (.A(n_11250_o_0),
    .B(n_11162_o_0),
    .Y(n_11580_o_0));
 OAI21xp33_ASAP7_75t_R n_11581 (.A1(n_11250_o_0),
    .A2(n_11162_o_0),
    .B(n_11580_o_0),
    .Y(n_11581_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11582 (.A1(n_11165_o_0),
    .A2(n_11581_o_0),
    .B(n_11559_o_0),
    .C(n_11202_o_0),
    .Y(n_11582_o_0));
 INVx1_ASAP7_75t_R n_11583 (.A(n_11520_o_0),
    .Y(n_11583_o_0));
 OAI21xp33_ASAP7_75t_R n_11584 (.A1(n_11192_o_0),
    .A2(n_11416_o_0),
    .B(n_11212_o_0),
    .Y(n_11584_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11585 (.A1(n_11583_o_0),
    .A2(n_11354_o_0),
    .B(n_11192_o_0),
    .C(n_11584_o_0),
    .Y(n_11585_o_0));
 AOI31xp33_ASAP7_75t_R n_11586 (.A1(n_11115_o_0),
    .A2(n_11579_o_0),
    .A3(n_11582_o_0),
    .B(n_11585_o_0),
    .Y(n_11586_o_0));
 AOI21xp33_ASAP7_75t_R n_11587 (.A1(n_11165_o_0),
    .A2(n_11448_o_0),
    .B(n_11208_o_0),
    .Y(n_11587_o_0));
 OAI21xp33_ASAP7_75t_R n_11588 (.A1(n_11190_o_0),
    .A2(n_11450_o_0),
    .B(n_11202_o_0),
    .Y(n_11588_o_0));
 INVx1_ASAP7_75t_R n_11589 (.A(n_11300_o_0),
    .Y(n_11589_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1159 (.A1(n_994_o_0),
    .A2(n_996_o_0),
    .B(n_878_o_0),
    .C(n_1028_o_0),
    .Y(n_1159_o_0));
 OAI22xp33_ASAP7_75t_R n_11590 (.A1(n_11587_o_0),
    .A2(n_11588_o_0),
    .B1(n_11275_o_0),
    .B2(n_11589_o_0),
    .Y(n_11590_o_0));
 OAI21xp33_ASAP7_75t_R n_11591 (.A1(net58),
    .A2(n_11190_o_0),
    .B(n_11250_o_0),
    .Y(n_11591_o_0));
 AOI21xp33_ASAP7_75t_R n_11592 (.A1(n_11239_o_0),
    .A2(n_11591_o_0),
    .B(n_11192_o_0),
    .Y(n_11592_o_0));
 NAND2xp33_ASAP7_75t_R n_11593 (.A(n_11239_o_0),
    .B(n_11192_o_0),
    .Y(n_11593_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11594 (.A1(n_11190_o_0),
    .A2(n_11137_o_0),
    .B(n_11334_o_0),
    .C(n_11593_o_0),
    .Y(n_11594_o_0));
 OAI21xp33_ASAP7_75t_R n_11595 (.A1(n_11592_o_0),
    .A2(n_11594_o_0),
    .B(n_11115_o_0),
    .Y(n_11595_o_0));
 OAI211xp5_ASAP7_75t_R n_11596 (.A1(n_11590_o_0),
    .A2(n_11115_o_0),
    .B(n_11393_o_0),
    .C(n_11595_o_0),
    .Y(n_11596_o_0));
 OAI21xp33_ASAP7_75t_R n_11597 (.A1(n_11106_o_0),
    .A2(n_11586_o_0),
    .B(n_11596_o_0),
    .Y(n_11597_o_0));
 AOI211xp5_ASAP7_75t_R n_11598 (.A1(n_11197_o_0),
    .A2(n_11454_o_0),
    .B(n_11397_o_0),
    .C(n_11266_o_0),
    .Y(n_11598_o_0));
 NAND3xp33_ASAP7_75t_R n_11599 (.A(n_11206_o_0),
    .B(n_11282_o_0),
    .C(n_11165_o_0),
    .Y(n_11599_o_0));
 OAI31xp33_ASAP7_75t_R n_1160 (.A1(net42),
    .A2(n_1159_o_0),
    .A3(n_1119_o_0),
    .B(n_904_o_0),
    .Y(n_1160_o_0));
 AOI21xp33_ASAP7_75t_R n_11600 (.A1(n_11205_o_0),
    .A2(n_11599_o_0),
    .B(n_11223_o_0),
    .Y(n_11600_o_0));
 OA21x2_ASAP7_75t_R n_11601 (.A1(n_11598_o_0),
    .A2(n_11600_o_0),
    .B(n_11192_o_0),
    .Y(n_11601_o_0));
 INVx1_ASAP7_75t_R n_11602 (.A(n_11466_o_0),
    .Y(n_11602_o_0));
 NOR2xp33_ASAP7_75t_R n_11603 (.A(n_11229_o_0),
    .B(n_11166_o_0),
    .Y(n_11603_o_0));
 AOI31xp33_ASAP7_75t_R n_11604 (.A1(n_11160_o_0),
    .A2(n_11243_o_0),
    .A3(n_11602_o_0),
    .B(n_11603_o_0),
    .Y(n_11604_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11605 (.A1(net35),
    .A2(net65),
    .B(n_11346_o_0),
    .C(n_11212_o_0),
    .Y(n_11605_o_0));
 OA21x2_ASAP7_75t_R n_11606 (.A1(n_11563_o_0),
    .A2(n_11251_o_0),
    .B(n_11605_o_0),
    .Y(n_11606_o_0));
 AOI211xp5_ASAP7_75t_R n_11607 (.A1(n_11604_o_0),
    .A2(n_11266_o_0),
    .B(net49),
    .C(n_11606_o_0),
    .Y(n_11607_o_0));
 OAI21xp33_ASAP7_75t_R n_11608 (.A1(n_11162_o_0),
    .A2(n_11197_o_0),
    .B(n_11554_o_0),
    .Y(n_11608_o_0));
 OAI31xp33_ASAP7_75t_R n_11609 (.A1(net37),
    .A2(n_11190_o_0),
    .A3(n_11162_o_0),
    .B(n_11608_o_0),
    .Y(n_11609_o_0));
 OAI221xp5_ASAP7_75t_R n_1161 (.A1(n_904_o_0),
    .A2(n_1154_o_0),
    .B1(n_1158_o_0),
    .B2(n_1160_o_0),
    .C(n_931_o_0),
    .Y(n_1161_o_0));
 NOR3xp33_ASAP7_75t_R n_11610 (.A(n_11160_o_0),
    .B(n_11186_o_0),
    .C(n_11152_o_0),
    .Y(n_11610_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11611 (.A1(n_11190_o_0),
    .A2(n_11189_o_0),
    .B(n_11223_o_0),
    .C(n_11610_o_0),
    .Y(n_11611_o_0));
 AOI21xp33_ASAP7_75t_R n_11612 (.A1(n_11160_o_0),
    .A2(n_11240_o_0),
    .B(n_11611_o_0),
    .Y(n_11612_o_0));
 AOI21xp33_ASAP7_75t_R n_11613 (.A1(n_11212_o_0),
    .A2(n_11609_o_0),
    .B(n_11612_o_0),
    .Y(n_11613_o_0));
 AOI21xp33_ASAP7_75t_R n_11614 (.A1(n_11327_o_0),
    .A2(n_11496_o_0),
    .B(n_11160_o_0),
    .Y(n_11614_o_0));
 INVx1_ASAP7_75t_R n_11615 (.A(n_11614_o_0),
    .Y(n_11615_o_0));
 OAI221xp5_ASAP7_75t_R n_11616 (.A1(n_11334_o_0),
    .A2(n_11465_o_0),
    .B1(n_11188_o_0),
    .B2(n_11231_o_0),
    .C(n_11615_o_0),
    .Y(n_11616_o_0));
 AOI21xp33_ASAP7_75t_R n_11617 (.A1(n_11250_o_0),
    .A2(n_11160_o_0),
    .B(n_11212_o_0),
    .Y(n_11617_o_0));
 NAND3xp33_ASAP7_75t_R n_11618 (.A(n_11496_o_0),
    .B(n_11282_o_0),
    .C(n_11165_o_0),
    .Y(n_11618_o_0));
 AOI21xp33_ASAP7_75t_R n_11619 (.A1(n_11617_o_0),
    .A2(n_11618_o_0),
    .B(n_11177_o_1),
    .Y(n_11619_o_0));
 OAI31xp33_ASAP7_75t_R n_1162 (.A1(n_931_o_0),
    .A2(n_1145_o_0),
    .A3(n_1151_o_0),
    .B(n_1161_o_0),
    .Y(n_1162_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11620 (.A1(n_11223_o_0),
    .A2(n_11616_o_0),
    .B(n_11619_o_0),
    .C(n_11105_o_0),
    .Y(n_11620_o_0));
 OAI21xp33_ASAP7_75t_R n_11621 (.A1(n_11202_o_0),
    .A2(n_11613_o_0),
    .B(n_11620_o_0),
    .Y(n_11621_o_0));
 OAI311xp33_ASAP7_75t_R n_11622 (.A1(n_11393_o_0),
    .A2(n_11601_o_0),
    .A3(n_11607_o_0),
    .B1(n_11221_o_0),
    .C1(n_11621_o_0),
    .Y(n_11622_o_0));
 OAI21xp33_ASAP7_75t_R n_11623 (.A1(n_11597_o_0),
    .A2(n_11221_o_0),
    .B(n_11622_o_0),
    .Y(n_11623_o_0));
 AOI31xp33_ASAP7_75t_R n_11624 (.A1(n_11162_o_0),
    .A2(n_11207_o_0),
    .A3(n_11196_o_0),
    .B(n_11200_o_0),
    .Y(n_11624_o_0));
 OAI211xp5_ASAP7_75t_R n_11625 (.A1(n_11162_o_0),
    .A2(n_11309_o_0),
    .B(n_11624_o_0),
    .C(n_11190_o_0),
    .Y(n_11625_o_0));
 OAI31xp33_ASAP7_75t_R n_11626 (.A1(net65),
    .A2(n_11624_o_0),
    .A3(n_11282_o_0),
    .B(n_11165_o_0),
    .Y(n_11626_o_0));
 AOI21xp33_ASAP7_75t_R n_11627 (.A1(n_11162_o_0),
    .A2(n_11309_o_0),
    .B(n_11160_o_0),
    .Y(n_11627_o_0));
 OR3x1_ASAP7_75t_R n_11628 (.A(n_11627_o_0),
    .B(n_11185_o_0),
    .C(net49),
    .Y(n_11628_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11629 (.A1(n_11625_o_0),
    .A2(n_11626_o_0),
    .B(n_11202_o_0),
    .C(n_11628_o_0),
    .Y(n_11629_o_0));
 NAND2xp33_ASAP7_75t_R n_1163 (.A(n_971_o_0),
    .B(n_1162_o_0),
    .Y(n_1163_o_0));
 NAND3xp33_ASAP7_75t_R n_11630 (.A(n_11580_o_0),
    .B(n_11179_o_0),
    .C(n_11190_o_0),
    .Y(n_11630_o_0));
 AOI22xp33_ASAP7_75t_R n_11631 (.A1(n_11259_o_0),
    .A2(n_11206_o_0),
    .B1(n_11160_o_0),
    .B2(net58),
    .Y(n_11631_o_0));
 OAI21xp33_ASAP7_75t_R n_11632 (.A1(n_11202_o_0),
    .A2(n_11631_o_0),
    .B(n_11223_o_0),
    .Y(n_11632_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11633 (.A1(n_11630_o_0),
    .A2(n_11380_o_0),
    .B(n_11632_o_0),
    .C(n_11105_o_0),
    .Y(n_11633_o_0));
 AOI211xp5_ASAP7_75t_R n_11634 (.A1(net58),
    .A2(net65),
    .B(n_11229_o_0),
    .C(n_11165_o_0),
    .Y(n_11634_o_0));
 NAND2xp33_ASAP7_75t_R n_11635 (.A(n_11450_o_0),
    .B(n_11185_o_0),
    .Y(n_11635_o_0));
 OAI211xp5_ASAP7_75t_R n_11636 (.A1(n_11387_o_0),
    .A2(n_11411_o_0),
    .B(n_11635_o_0),
    .C(n_11212_o_0),
    .Y(n_11636_o_0));
 OAI31xp33_ASAP7_75t_R n_11637 (.A1(n_11339_o_0),
    .A2(n_11614_o_0),
    .A3(n_11634_o_0),
    .B(n_11636_o_0),
    .Y(n_11637_o_0));
 AOI21xp33_ASAP7_75t_R n_11638 (.A1(n_11520_o_0),
    .A2(n_11334_o_0),
    .B(n_11266_o_0),
    .Y(n_11638_o_0));
 NAND2xp33_ASAP7_75t_R n_11639 (.A(n_11496_o_0),
    .B(n_11259_o_0),
    .Y(n_11639_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1164 (.A1(n_1130_o_0),
    .A2(n_1139_o_0),
    .B(n_971_o_0),
    .C(n_1163_o_0),
    .Y(n_1164_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11640 (.A1(n_11465_o_0),
    .A2(n_11334_o_0),
    .B(n_11639_o_0),
    .C(n_11115_o_0),
    .Y(n_11640_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11641 (.A1(n_11638_o_0),
    .A2(n_11640_o_0),
    .B(n_11202_o_0),
    .C(n_11296_o_0),
    .Y(n_11641_o_0));
 OAI21xp33_ASAP7_75t_R n_11642 (.A1(n_11224_o_0),
    .A2(n_11637_o_0),
    .B(n_11641_o_0),
    .Y(n_11642_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11643 (.A1(n_11266_o_0),
    .A2(n_11629_o_0),
    .B(n_11633_o_0),
    .C(n_11642_o_0),
    .Y(n_11643_o_0));
 AOI21xp33_ASAP7_75t_R n_11644 (.A1(n_11442_o_0),
    .A2(n_11198_o_0),
    .B(n_11192_o_0),
    .Y(n_11644_o_0));
 NAND4xp25_ASAP7_75t_R n_11645 (.A(n_11201_o_0),
    .B(n_11503_o_0),
    .C(n_11450_o_0),
    .D(n_11190_o_0),
    .Y(n_11645_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11646 (.A1(net58),
    .A2(net65),
    .B(n_11250_o_0),
    .C(n_11160_o_0),
    .Y(n_11646_o_0));
 OAI31xp33_ASAP7_75t_R n_11647 (.A1(n_11190_o_0),
    .A2(n_11465_o_0),
    .A3(n_11466_o_0),
    .B(n_11646_o_0),
    .Y(n_11647_o_0));
 AOI22xp33_ASAP7_75t_R n_11648 (.A1(n_11644_o_0),
    .A2(n_11645_o_0),
    .B1(n_11192_o_0),
    .B2(n_11647_o_0),
    .Y(n_11648_o_0));
 NAND3xp33_ASAP7_75t_R n_11649 (.A(n_11618_o_0),
    .B(n_11317_o_0),
    .C(n_11177_o_1),
    .Y(n_11649_o_0));
 AND4x1_ASAP7_75t_R n_1165 (.A(n_1045_o_0),
    .B(n_1085_o_0),
    .C(n_985_o_0),
    .D(net16),
    .Y(n_1165_o_0));
 OAI31xp33_ASAP7_75t_R n_11650 (.A1(n_11188_o_0),
    .A2(n_11165_o_0),
    .A3(n_11162_o_0),
    .B(n_11224_o_0),
    .Y(n_11650_o_0));
 AOI31xp33_ASAP7_75t_R n_11651 (.A1(n_11250_o_0),
    .A2(net65),
    .A3(n_11165_o_0),
    .B(n_11650_o_0),
    .Y(n_11651_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11652 (.A1(n_11250_o_0),
    .A2(net58),
    .B(net65),
    .C(n_11651_o_0),
    .Y(n_11652_o_0));
 AOI21xp33_ASAP7_75t_R n_11653 (.A1(n_11649_o_0),
    .A2(n_11652_o_0),
    .B(n_11115_o_0),
    .Y(n_11653_o_0));
 AOI211xp5_ASAP7_75t_R n_11654 (.A1(n_11223_o_0),
    .A2(n_11648_o_0),
    .B(n_11653_o_0),
    .C(n_11296_o_0),
    .Y(n_11654_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11655 (.A1(net35),
    .A2(n_11162_o_0),
    .B(n_11165_o_0),
    .C(n_11430_o_0),
    .Y(n_11655_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11656 (.A1(n_11454_o_0),
    .A2(n_11187_o_0),
    .B(n_11655_o_0),
    .C(n_11202_o_0),
    .Y(n_11656_o_0));
 OAI21xp33_ASAP7_75t_R n_11657 (.A1(net65),
    .A2(n_11197_o_0),
    .B(n_11209_o_0),
    .Y(n_11657_o_0));
 OAI21xp33_ASAP7_75t_R n_11658 (.A1(n_11314_o_0),
    .A2(n_11281_o_0),
    .B(n_11657_o_0),
    .Y(n_11658_o_0));
 AOI21xp33_ASAP7_75t_R n_11659 (.A1(n_11192_o_0),
    .A2(n_11658_o_0),
    .B(n_11115_o_0),
    .Y(n_11659_o_0));
 INVx1_ASAP7_75t_R n_1166 (.A(n_1004_o_0),
    .Y(n_1166_o_0));
 NAND3xp33_ASAP7_75t_R n_11660 (.A(n_11206_o_0),
    .B(n_11282_o_0),
    .C(n_11160_o_0),
    .Y(n_11660_o_0));
 NAND3xp33_ASAP7_75t_R n_11661 (.A(n_11660_o_0),
    .B(n_11343_o_0),
    .C(n_11177_o_1),
    .Y(n_11661_o_0));
 AO21x1_ASAP7_75t_R n_11662 (.A1(n_11165_o_0),
    .A2(n_11291_o_0),
    .B(n_11650_o_0),
    .Y(n_11662_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11663 (.A1(n_11661_o_0),
    .A2(n_11662_o_0),
    .B(n_11212_o_0),
    .C(n_11105_o_0),
    .Y(n_11663_o_0));
 AOI21xp33_ASAP7_75t_R n_11664 (.A1(n_11656_o_0),
    .A2(n_11659_o_0),
    .B(n_11663_o_0),
    .Y(n_11664_o_0));
 OAI21xp33_ASAP7_75t_R n_11665 (.A1(n_11654_o_0),
    .A2(n_11664_o_0),
    .B(n_11221_o_0),
    .Y(n_11665_o_0));
 OAI21xp33_ASAP7_75t_R n_11666 (.A1(n_11221_o_0),
    .A2(n_11643_o_0),
    .B(n_11665_o_0),
    .Y(n_11666_o_0));
 INVx1_ASAP7_75t_R n_11667 (.A(_00962_),
    .Y(n_11667_o_0));
 XOR2xp5_ASAP7_75t_R n_11668 (.A(_01025_),
    .B(_01112_),
    .Y(n_11668_o_0));
 XNOR2xp5_ASAP7_75t_R n_11669 (.A(_01026_),
    .B(n_11668_o_0),
    .Y(n_11669_o_0));
 OAI21xp33_ASAP7_75t_R n_1167 (.A1(n_836_o_0),
    .A2(n_913_o_0),
    .B(n_877_o_0),
    .Y(n_1167_o_0));
 NAND2xp33_ASAP7_75t_R n_11670 (.A(n_4824_o_0),
    .B(n_11669_o_0),
    .Y(n_11670_o_0));
 OAI21xp33_ASAP7_75t_R n_11671 (.A1(n_4824_o_0),
    .A2(n_11669_o_0),
    .B(n_11670_o_0),
    .Y(n_11671_o_0));
 NOR2xp33_ASAP7_75t_R n_11672 (.A(_00725_),
    .B(net),
    .Y(n_11672_o_0));
 AOI21xp33_ASAP7_75t_R n_11673 (.A1(net),
    .A2(n_11671_o_0),
    .B(n_11672_o_0),
    .Y(n_11673_o_0));
 HAxp5_ASAP7_75t_R n_11674 (.A(n_11667_o_0),
    .B(n_11673_o_0),
    .CON(n_11674_o_0),
    .SN(n_11674_o_1));
 INVx1_ASAP7_75t_R n_11675 (.A(n_11674_o_1),
    .Y(n_11675_o_0));
 XNOR2xp5_ASAP7_75t_R n_11676 (.A(_01026_),
    .B(_01113_),
    .Y(n_11676_o_0));
 XNOR2xp5_ASAP7_75t_R n_11677 (.A(n_4887_o_0),
    .B(n_11676_o_0),
    .Y(n_11677_o_0));
 NOR2xp33_ASAP7_75t_R n_11678 (.A(n_4813_o_0),
    .B(n_11677_o_0),
    .Y(n_11678_o_0));
 NOR2xp33_ASAP7_75t_R n_11679 (.A(_00724_),
    .B(net),
    .Y(n_11679_o_0));
 OAI21xp33_ASAP7_75t_R n_1168 (.A1(n_892_o_0),
    .A2(n_1167_o_0),
    .B(n_891_o_0),
    .Y(n_1168_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11680 (.A1(n_4813_o_0),
    .A2(n_11677_o_0),
    .B(n_11678_o_0),
    .C(net),
    .D(n_11679_o_0),
    .Y(n_11680_o_0));
 HAxp5_ASAP7_75t_R n_11681 (.A(n_11680_o_0),
    .B(n_1858_o_0),
    .CON(n_11681_o_0),
    .SN(n_11681_o_1));
 XNOR2xp5_ASAP7_75t_R n_11682 (.A(_01033_),
    .B(_01073_),
    .Y(n_11682_o_0));
 XNOR2xp5_ASAP7_75t_R n_11683 (.A(_01111_),
    .B(n_11682_o_0),
    .Y(n_11683_o_0));
 XOR2xp5_ASAP7_75t_R n_11684 (.A(_01024_),
    .B(_01025_),
    .Y(n_11684_o_0));
 NOR2xp33_ASAP7_75t_R n_11685 (.A(n_11684_o_0),
    .B(n_11683_o_0),
    .Y(n_11685_o_0));
 NOR2xp33_ASAP7_75t_R n_11686 (.A(_00726_),
    .B(net),
    .Y(n_11686_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11687 (.A1(n_11683_o_0),
    .A2(n_11684_o_0),
    .B(n_11685_o_0),
    .C(net39),
    .D(n_11686_o_0),
    .Y(n_11687_o_0));
 XNOR2xp5_ASAP7_75t_R n_11688 (.A(_00961_),
    .B(n_11687_o_0),
    .Y(n_11688_o_0));
 INVx1_ASAP7_75t_R n_11689 (.A(n_11688_o_0),
    .Y(n_11689_o_0));
 AOI21xp33_ASAP7_75t_R n_1169 (.A1(n_1166_o_0),
    .A2(n_1005_o_0),
    .B(n_1168_o_0),
    .Y(n_1169_o_0));
 NAND2xp33_ASAP7_75t_R n_11690 (.A(n_9446_o_0),
    .B(n_4862_o_0),
    .Y(n_11690_o_0));
 XNOR2xp5_ASAP7_75t_R n_11691 (.A(_01069_),
    .B(n_4900_o_0),
    .Y(n_11691_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11692 (.A1(_01107_),
    .A2(_01114_),
    .B(n_9445_o_0),
    .C(n_4861_o_0),
    .Y(n_11692_o_0));
 AOI31xp33_ASAP7_75t_R n_11693 (.A1(n_11690_o_0),
    .A2(n_11691_o_0),
    .A3(n_11692_o_0),
    .B(n_3021_o_0),
    .Y(n_11693_o_0));
 NOR2xp33_ASAP7_75t_R n_11694 (.A(_01069_),
    .B(n_4915_o_0),
    .Y(n_11694_o_0));
 INVx1_ASAP7_75t_R n_11695 (.A(_01069_),
    .Y(n_11695_o_0));
 NOR2xp33_ASAP7_75t_R n_11696 (.A(n_11695_o_0),
    .B(n_4900_o_0),
    .Y(n_11696_o_0));
 OAI21xp33_ASAP7_75t_R n_11697 (.A1(n_4861_o_0),
    .A2(n_9437_o_0),
    .B(n_11692_o_0),
    .Y(n_11697_o_0));
 OAI21xp33_ASAP7_75t_R n_11698 (.A1(n_11694_o_0),
    .A2(n_11696_o_0),
    .B(n_11697_o_0),
    .Y(n_11698_o_0));
 AOI22xp33_ASAP7_75t_R n_11699 (.A1(n_11693_o_0),
    .A2(n_11698_o_0),
    .B1(net3),
    .B2(_00410_),
    .Y(n_11699_o_0));
 NAND2xp33_ASAP7_75t_R n_1170 (.A(n_956_o_0),
    .B(n_1166_o_0),
    .Y(n_1170_o_0));
 INVx1_ASAP7_75t_R n_11700 (.A(_00957_),
    .Y(n_11700_o_0));
 INVx1_ASAP7_75t_R n_11701 (.A(_00410_),
    .Y(n_11701_o_0));
 NAND2xp33_ASAP7_75t_R n_11702 (.A(n_11695_o_0),
    .B(n_4900_o_0),
    .Y(n_11702_o_0));
 OAI21xp33_ASAP7_75t_R n_11703 (.A1(n_4900_o_0),
    .A2(n_11695_o_0),
    .B(n_11702_o_0),
    .Y(n_11703_o_0));
 OAI21xp33_ASAP7_75t_R n_11704 (.A1(n_11697_o_0),
    .A2(n_11703_o_0),
    .B(net39),
    .Y(n_11704_o_0));
 INVx1_ASAP7_75t_R n_11705 (.A(n_11698_o_0),
    .Y(n_11705_o_0));
 OAI221xp5_ASAP7_75t_R n_11706 (.A1(net39),
    .A2(n_11701_o_0),
    .B1(n_11704_o_0),
    .B2(n_11705_o_0),
    .C(n_11700_o_0),
    .Y(n_11706_o_0));
 OAI21x1_ASAP7_75t_R n_11707 (.A1(n_11699_o_0),
    .A2(n_11700_o_0),
    .B(n_11706_o_0),
    .Y(n_11707_o_0));
 NAND2xp33_ASAP7_75t_R n_11708 (.A(n_4884_o_0),
    .B(n_4915_o_0),
    .Y(n_11708_o_0));
 OAI21xp33_ASAP7_75t_R n_11709 (.A1(n_4915_o_0),
    .A2(n_4884_o_0),
    .B(n_11708_o_0),
    .Y(n_11709_o_0));
 OAI31xp33_ASAP7_75t_R n_1171 (.A1(n_878_o_0),
    .A2(n_1025_o_0),
    .A3(n_938_o_0),
    .B(n_1170_o_0),
    .Y(n_1171_o_0));
 NOR2xp33_ASAP7_75t_R n_11710 (.A(n_4900_o_0),
    .B(n_4891_o_0),
    .Y(n_11710_o_0));
 AOI211xp5_ASAP7_75t_R n_11711 (.A1(n_4900_o_0),
    .A2(n_4891_o_0),
    .B(n_11710_o_0),
    .C(_01114_),
    .Y(n_11711_o_0));
 NOR2xp33_ASAP7_75t_R n_11712 (.A(_00411_),
    .B(_00858_),
    .Y(n_11712_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11713 (.A1(n_11709_o_0),
    .A2(_01114_),
    .B(n_11711_o_0),
    .C(net77),
    .D(n_11712_o_0),
    .Y(n_11713_o_0));
 INVx1_ASAP7_75t_R n_11714 (.A(_01114_),
    .Y(n_11714_o_0));
 OAI211xp5_ASAP7_75t_R n_11715 (.A1(n_4915_o_0),
    .A2(n_4884_o_0),
    .B(n_11708_o_0),
    .C(n_11714_o_0),
    .Y(n_11715_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11716 (.A1(n_4900_o_0),
    .A2(n_4891_o_0),
    .B(n_11710_o_0),
    .C(_01114_),
    .Y(n_11716_o_0));
 INVx1_ASAP7_75t_R n_11717 (.A(n_11712_o_0),
    .Y(n_11717_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11718 (.A1(n_11715_o_0),
    .A2(n_11716_o_0),
    .B(net1),
    .C(n_11717_o_0),
    .D(_00956_),
    .Y(n_11718_o_0));
 AO21x1_ASAP7_75t_R n_11719 (.A1(_00956_),
    .A2(n_11713_o_0),
    .B(n_11718_o_0),
    .Y(n_11719_o_0));
 OAI21xp33_ASAP7_75t_R n_1172 (.A1(n_887_o_0),
    .A2(n_996_o_0),
    .B(n_878_o_0),
    .Y(n_1172_o_0));
 INVx1_ASAP7_75t_R n_11720 (.A(_00958_),
    .Y(n_11720_o_0));
 XNOR2xp5_ASAP7_75t_R n_11721 (.A(_01021_),
    .B(_01108_),
    .Y(n_11721_o_0));
 NAND2xp33_ASAP7_75t_R n_11722 (.A(n_4865_o_0),
    .B(n_11721_o_0),
    .Y(n_11722_o_0));
 OAI21xp33_ASAP7_75t_R n_11723 (.A1(n_11721_o_0),
    .A2(n_4865_o_0),
    .B(n_11722_o_0),
    .Y(n_11723_o_0));
 NOR2xp33_ASAP7_75t_R n_11724 (.A(n_4865_o_0),
    .B(n_11721_o_0),
    .Y(n_11724_o_0));
 AOI211xp5_ASAP7_75t_R n_11725 (.A1(n_11721_o_0),
    .A2(n_4865_o_0),
    .B(n_11724_o_0),
    .C(n_9424_o_0),
    .Y(n_11725_o_0));
 NOR2xp33_ASAP7_75t_R n_11726 (.A(_00413_),
    .B(_00858_),
    .Y(n_11726_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11727 (.A1(n_9424_o_0),
    .A2(n_11723_o_0),
    .B(n_11725_o_0),
    .C(net77),
    .D(n_11726_o_0),
    .Y(n_11727_o_0));
 INVx1_ASAP7_75t_R n_11728 (.A(n_9424_o_0),
    .Y(n_11728_o_0));
 OAI211xp5_ASAP7_75t_R n_11729 (.A1(n_11721_o_0),
    .A2(n_4865_o_0),
    .B(n_11722_o_0),
    .C(n_11728_o_0),
    .Y(n_11729_o_0));
 NAND4xp25_ASAP7_75t_R n_1173 (.A(n_1172_o_0),
    .B(n_1002_o_0),
    .C(n_985_o_0),
    .D(n_891_o_0),
    .Y(n_1173_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11730 (.A1(n_11721_o_0),
    .A2(n_4865_o_0),
    .B(n_11724_o_0),
    .C(n_9424_o_0),
    .Y(n_11730_o_0));
 INVx1_ASAP7_75t_R n_11731 (.A(n_11726_o_0),
    .Y(n_11731_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11732 (.A1(n_11729_o_0),
    .A2(n_11730_o_0),
    .B(net3),
    .C(n_11731_o_0),
    .D(n_11720_o_0),
    .Y(n_11732_o_0));
 AOI21x1_ASAP7_75t_R n_11733 (.A1(n_11720_o_0),
    .A2(n_11727_o_0),
    .B(n_11732_o_0),
    .Y(n_11733_o_0));
 XNOR2xp5_ASAP7_75t_R n_11734 (.A(_01071_),
    .B(n_4834_o_0),
    .Y(n_11734_o_0));
 OAI211xp5_ASAP7_75t_R n_11735 (.A1(n_9455_o_0),
    .A2(n_9456_o_0),
    .B(n_11734_o_0),
    .C(n_9457_o_0),
    .Y(n_11735_o_0));
 NOR2xp33_ASAP7_75t_R n_11736 (.A(_01071_),
    .B(n_4839_o_0),
    .Y(n_11736_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11737 (.A1(_01071_),
    .A2(n_4839_o_0),
    .B(n_11736_o_0),
    .C(n_9458_o_0),
    .Y(n_11737_o_0));
 NOR2xp33_ASAP7_75t_R n_11738 (.A(_00728_),
    .B(_00858_),
    .Y(n_11738_o_0));
 INVx1_ASAP7_75t_R n_11739 (.A(n_11738_o_0),
    .Y(n_11739_o_0));
 OAI211xp5_ASAP7_75t_R n_1174 (.A1(n_1171_o_0),
    .A2(net14),
    .B(n_1173_o_0),
    .C(n_903_o_0),
    .Y(n_1174_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11740 (.A1(n_11735_o_0),
    .A2(n_11737_o_0),
    .B(net5),
    .C(n_11739_o_0),
    .Y(n_11740_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11741 (.A1(n_11737_o_0),
    .A2(n_11735_o_0),
    .B(net9),
    .C(n_11739_o_0),
    .D(_00959_),
    .Y(n_11741_o_0));
 INVx1_ASAP7_75t_R n_11742 (.A(n_11741_o_0),
    .Y(n_11742_o_0));
 OAI21x1_ASAP7_75t_R n_11743 (.A1(n_1922_o_0),
    .A2(n_11740_o_0),
    .B(n_11742_o_0),
    .Y(n_11743_o_0));
 OAI21xp33_ASAP7_75t_R n_11744 (.A1(n_11733_o_0),
    .A2(n_11719_o_0),
    .B(n_11743_o_0),
    .Y(n_11744_o_0));
 AOI21xp33_ASAP7_75t_R n_11745 (.A1(n_11707_o_0),
    .A2(n_11719_o_0),
    .B(n_11744_o_0),
    .Y(n_11745_o_0));
 AOI21xp33_ASAP7_75t_R n_11746 (.A1(n_11697_o_0),
    .A2(n_11703_o_0),
    .B(n_11704_o_0),
    .Y(n_11746_o_0));
 AOI221xp5_ASAP7_75t_R n_11747 (.A1(net1),
    .A2(_00410_),
    .B1(n_11698_o_0),
    .B2(n_11693_o_0),
    .C(_00957_),
    .Y(n_11747_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11748 (.A1(net9),
    .A2(_00410_),
    .B(n_11746_o_0),
    .C(_00957_),
    .D(n_11747_o_0),
    .Y(n_11748_o_0));
 HAxp5_ASAP7_75t_R n_11749 (.A(n_11719_o_0),
    .B(n_11748_o_0),
    .CON(n_11749_o_0),
    .SN(n_11749_o_1));
 OAI31xp33_ASAP7_75t_R n_1175 (.A1(n_1165_o_0),
    .A2(n_1169_o_0),
    .A3(n_903_o_0),
    .B(n_1174_o_0),
    .Y(n_1175_o_0));
 NAND2xp33_ASAP7_75t_R n_11750 (.A(_00959_),
    .B(n_11740_o_0),
    .Y(n_11750_o_0));
 OAI21x1_ASAP7_75t_R n_11751 (.A1(_00959_),
    .A2(n_11740_o_0),
    .B(n_11750_o_0),
    .Y(n_11751_o_0));
 AOI21xp5_ASAP7_75t_R n_11752 (.A1(_00956_),
    .A2(n_11713_o_0),
    .B(n_11718_o_0),
    .Y(n_11752_o_0));
 NAND2xp33_ASAP7_75t_R n_11753 (.A(n_11733_o_0),
    .B(n_11752_o_0),
    .Y(n_11753_o_0));
 NAND3xp33_ASAP7_75t_R n_11754 (.A(n_11749_o_0),
    .B(n_11751_o_0),
    .C(n_11753_o_0),
    .Y(n_11754_o_0));
 INVx1_ASAP7_75t_R n_11755 (.A(n_11754_o_0),
    .Y(n_11755_o_0));
 XNOR2xp5_ASAP7_75t_R n_11756 (.A(_01072_),
    .B(n_4961_o_0),
    .Y(n_11756_o_0));
 XOR2xp5_ASAP7_75t_R n_11757 (.A(n_11756_o_0),
    .B(n_9496_o_0),
    .Y(n_11757_o_0));
 NOR2xp33_ASAP7_75t_R n_11758 (.A(_00727_),
    .B(net39),
    .Y(n_11758_o_0));
 AOI21xp33_ASAP7_75t_R n_11759 (.A1(net),
    .A2(n_11757_o_0),
    .B(n_11758_o_0),
    .Y(n_11759_o_0));
 AOI21xp33_ASAP7_75t_R n_1176 (.A1(n_956_o_0),
    .A2(n_910_o_0),
    .B(n_877_o_0),
    .Y(n_1176_o_0));
 NAND2xp33_ASAP7_75t_R n_11760 (.A(_00960_),
    .B(n_11759_o_0),
    .Y(n_11760_o_0));
 OAI21xp5_ASAP7_75t_R n_11761 (.A1(_00960_),
    .A2(n_11759_o_0),
    .B(n_11760_o_0),
    .Y(n_11761_o_0));
 NOR2xp33_ASAP7_75t_R n_11762 (.A(_00959_),
    .B(n_11740_o_0),
    .Y(n_11762_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11763 (.A1(n_11740_o_0),
    .A2(_00959_),
    .B(n_11762_o_0),
    .C(n_11733_o_0),
    .Y(n_11763_o_0));
 NOR2xp67_ASAP7_75t_R n_11764 (.A(n_11752_o_0),
    .B(n_11748_o_0),
    .Y(n_11764_o_0));
 NOR2xp33_ASAP7_75t_R n_11765 (.A(n_11707_o_0),
    .B(n_11753_o_0),
    .Y(n_11765_o_0));
 AO21x1_ASAP7_75t_R n_11766 (.A1(n_11720_o_0),
    .A2(n_11727_o_0),
    .B(n_11732_o_0),
    .Y(n_11766_o_0));
 NAND2xp33_ASAP7_75t_R n_11767 (.A(n_11752_o_0),
    .B(n_11707_o_0),
    .Y(n_11767_o_0));
 OAI311xp33_ASAP7_75t_R n_11768 (.A1(n_11694_o_0),
    .A2(n_11696_o_0),
    .A3(n_11697_o_0),
    .B1(net),
    .C1(n_11698_o_0),
    .Y(n_11768_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11769 (.A1(n_11701_o_0),
    .A2(net),
    .B(n_11768_o_0),
    .C(n_11700_o_0),
    .Y(n_11769_o_0));
 OA21x2_ASAP7_75t_R n_1177 (.A1(n_1057_o_0),
    .A2(n_1176_o_0),
    .B(net14),
    .Y(n_1177_o_0));
 AOI21xp33_ASAP7_75t_R n_11770 (.A1(n_11715_o_0),
    .A2(n_11716_o_0),
    .B(net2),
    .Y(n_11770_o_0));
 INVx1_ASAP7_75t_R n_11771 (.A(_00956_),
    .Y(n_11771_o_0));
 AOI211xp5_ASAP7_75t_R n_11772 (.A1(n_11712_o_0),
    .A2(net2),
    .B(n_11770_o_0),
    .C(n_11771_o_0),
    .Y(n_11772_o_0));
 OAI22xp33_ASAP7_75t_R n_11773 (.A1(n_11747_o_0),
    .A2(n_11769_o_0),
    .B1(n_11772_o_0),
    .B2(n_11718_o_0),
    .Y(n_11773_o_0));
 OAI21xp5_ASAP7_75t_R n_11774 (.A1(n_11707_o_0),
    .A2(n_11719_o_0),
    .B(n_11773_o_0),
    .Y(n_11774_o_0));
 INVx1_ASAP7_75t_R n_11775 (.A(n_11734_o_0),
    .Y(n_11775_o_0));
 OAI21xp33_ASAP7_75t_R n_11776 (.A1(n_9458_o_0),
    .A2(n_11775_o_0),
    .B(n_11737_o_0),
    .Y(n_11776_o_0));
 AOI211xp5_ASAP7_75t_R n_11777 (.A1(n_11776_o_0),
    .A2(net39),
    .B(n_1922_o_0),
    .C(n_11738_o_0),
    .Y(n_11777_o_0));
 NOR2xp67_ASAP7_75t_R n_11778 (.A(n_11741_o_0),
    .B(n_11777_o_0),
    .Y(n_11778_o_0));
 AOI21xp33_ASAP7_75t_R n_11779 (.A1(n_11766_o_0),
    .A2(n_11774_o_0),
    .B(n_11778_o_0),
    .Y(n_11779_o_0));
 AOI22xp33_ASAP7_75t_R n_1178 (.A1(n_860_o_0),
    .A2(n_881_o_0),
    .B1(n_1005_o_0),
    .B2(n_878_o_0),
    .Y(n_1178_o_0));
 AOI31xp33_ASAP7_75t_R n_11780 (.A1(n_11766_o_0),
    .A2(n_11751_o_0),
    .A3(n_11767_o_0),
    .B(n_11779_o_0),
    .Y(n_11780_o_0));
 AOI211xp5_ASAP7_75t_R n_11781 (.A1(n_11757_o_0),
    .A2(net),
    .B(_00960_),
    .C(n_11758_o_0),
    .Y(n_11781_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_11782 (.A1(n_11757_o_0),
    .A2(net),
    .B(n_11758_o_0),
    .C(_00960_),
    .D(n_11781_o_0),
    .Y(n_11782_o_0));
 OAI221xp5_ASAP7_75t_R n_11783 (.A1(n_11763_o_0),
    .A2(n_11764_o_0),
    .B1(n_11765_o_0),
    .B2(n_11780_o_0),
    .C(n_11782_o_0),
    .Y(n_11783_o_0));
 OAI31xp33_ASAP7_75t_R n_11784 (.A1(n_11745_o_0),
    .A2(n_11755_o_0),
    .A3(n_11761_o_0),
    .B(n_11783_o_0),
    .Y(n_11784_o_0));
 INVx1_ASAP7_75t_R n_11785 (.A(n_11774_o_0),
    .Y(n_11785_o_0));
 OAI21xp33_ASAP7_75t_R n_11786 (.A1(n_11733_o_0),
    .A2(n_11785_o_0),
    .B(n_11778_o_0),
    .Y(n_11786_o_0));
 AOI21xp33_ASAP7_75t_R n_11787 (.A1(n_11752_o_0),
    .A2(n_11707_o_0),
    .B(n_11766_o_0),
    .Y(n_11787_o_0));
 NOR2xp33_ASAP7_75t_R n_11788 (.A(n_11733_o_0),
    .B(n_11764_o_0),
    .Y(n_11788_o_0));
 AOI21xp5_ASAP7_75t_R n_11789 (.A1(n_11740_o_0),
    .A2(_00959_),
    .B(n_11762_o_0),
    .Y(n_11789_o_0));
 OAI21xp33_ASAP7_75t_R n_1179 (.A1(n_1178_o_0),
    .A2(net14),
    .B(n_904_o_0),
    .Y(n_1179_o_0));
 OAI21xp33_ASAP7_75t_R n_11790 (.A1(n_11787_o_0),
    .A2(n_11788_o_0),
    .B(n_11789_o_0),
    .Y(n_11790_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11791 (.A1(n_11733_o_0),
    .A2(n_11764_o_0),
    .B(n_11786_o_0),
    .C(n_11790_o_0),
    .Y(n_11791_o_0));
 NOR2xp33_ASAP7_75t_R n_11792 (.A(n_11766_o_0),
    .B(n_11707_o_0),
    .Y(n_11792_o_0));
 INVx1_ASAP7_75t_R n_11793 (.A(n_11792_o_0),
    .Y(n_11793_o_0));
 OAI21xp33_ASAP7_75t_R n_11794 (.A1(n_11733_o_0),
    .A2(n_11774_o_0),
    .B(n_11743_o_0),
    .Y(n_11794_o_0));
 INVx1_ASAP7_75t_R n_11795 (.A(n_11794_o_0),
    .Y(n_11795_o_0));
 INVx1_ASAP7_75t_R n_11796 (.A(n_11761_o_0),
    .Y(n_11796_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11797 (.A1(n_11774_o_0),
    .A2(n_11733_o_0),
    .B(n_11789_o_0),
    .C(n_11796_o_0),
    .Y(n_11797_o_0));
 XNOR2xp5_ASAP7_75t_R n_11798 (.A(n_1877_o_0),
    .B(n_11687_o_0),
    .Y(n_11798_o_0));
 INVx1_ASAP7_75t_R n_11799 (.A(n_11798_o_0),
    .Y(n_11799_o_0));
 NOR2xp33_ASAP7_75t_R n_1180 (.A(n_989_o_0),
    .B(n_915_o_0),
    .Y(n_1180_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11800 (.A1(n_11793_o_0),
    .A2(n_11795_o_0),
    .B(n_11797_o_0),
    .C(n_11799_o_0),
    .Y(n_11800_o_0));
 AOI21xp33_ASAP7_75t_R n_11801 (.A1(n_11782_o_0),
    .A2(n_11791_o_0),
    .B(n_11800_o_0),
    .Y(n_11801_o_0));
 AOI21xp33_ASAP7_75t_R n_11802 (.A1(n_11689_o_0),
    .A2(n_11784_o_0),
    .B(n_11801_o_0),
    .Y(n_11802_o_0));
 INVx1_ASAP7_75t_R n_11803 (.A(n_11767_o_0),
    .Y(n_11803_o_0));
 OAI21xp33_ASAP7_75t_R n_11804 (.A1(n_11766_o_0),
    .A2(n_11803_o_0),
    .B(n_11778_o_0),
    .Y(n_11804_o_0));
 NAND2xp33_ASAP7_75t_R n_11805 (.A(n_11766_o_0),
    .B(n_11719_o_0),
    .Y(n_11805_o_0));
 NOR2xp33_ASAP7_75t_R n_11806 (.A(n_11707_o_0),
    .B(n_11805_o_0),
    .Y(n_11806_o_0));
 NAND2xp33_ASAP7_75t_R n_11807 (.A(n_11766_o_0),
    .B(n_11764_o_0),
    .Y(n_11807_o_0));
 OAI22xp33_ASAP7_75t_R n_11808 (.A1(n_11804_o_0),
    .A2(n_11806_o_0),
    .B1(n_11807_o_0),
    .B2(n_11751_o_0),
    .Y(n_11808_o_0));
 NAND3xp33_ASAP7_75t_R n_11809 (.A(n_11707_o_0),
    .B(n_11752_o_0),
    .C(n_11733_o_0),
    .Y(n_11809_o_0));
 OAI21xp33_ASAP7_75t_R n_1181 (.A1(n_847_o_0),
    .A2(n_859_o_0),
    .B(n_953_o_0),
    .Y(n_1181_o_0));
 NAND2xp33_ASAP7_75t_R n_11810 (.A(n_11743_o_0),
    .B(n_11809_o_0),
    .Y(n_11810_o_0));
 NAND2xp33_ASAP7_75t_R n_11811 (.A(n_11766_o_0),
    .B(n_11719_o_0),
    .Y(n_11811_o_0));
 NOR2xp33_ASAP7_75t_R n_11812 (.A(n_11707_o_0),
    .B(n_11811_o_0),
    .Y(n_11812_o_0));
 NAND3xp33_ASAP7_75t_R n_11813 (.A(n_11764_o_0),
    .B(n_11751_o_0),
    .C(n_11766_o_0),
    .Y(n_11813_o_0));
 OAI211xp5_ASAP7_75t_R n_11814 (.A1(n_11810_o_0),
    .A2(n_11812_o_0),
    .B(n_11813_o_0),
    .C(n_11796_o_0),
    .Y(n_11814_o_0));
 OAI21xp33_ASAP7_75t_R n_11815 (.A1(n_11796_o_0),
    .A2(n_11808_o_0),
    .B(n_11814_o_0),
    .Y(n_11815_o_0));
 NAND2xp33_ASAP7_75t_R n_11816 (.A(n_11719_o_0),
    .B(n_11748_o_0),
    .Y(n_11816_o_0));
 NAND2xp33_ASAP7_75t_R n_11817 (.A(n_11733_o_0),
    .B(n_11816_o_0),
    .Y(n_11817_o_0));
 OAI211xp5_ASAP7_75t_R n_11818 (.A1(n_11707_o_0),
    .A2(n_11805_o_0),
    .B(n_11817_o_0),
    .C(n_11789_o_0),
    .Y(n_11818_o_0));
 NAND2xp33_ASAP7_75t_R n_11819 (.A(n_11733_o_0),
    .B(n_11764_o_0),
    .Y(n_11819_o_0));
 AOI21xp33_ASAP7_75t_R n_1182 (.A1(n_877_o_0),
    .A2(n_1181_o_0),
    .B(n_891_o_0),
    .Y(n_1182_o_0));
 INVx1_ASAP7_75t_R n_11820 (.A(n_11753_o_0),
    .Y(n_11820_o_0));
 OAI31xp33_ASAP7_75t_R n_11821 (.A1(n_11733_o_0),
    .A2(n_11764_o_0),
    .A3(n_11743_o_0),
    .B(n_11761_o_0),
    .Y(n_11821_o_0));
 AOI21xp33_ASAP7_75t_R n_11822 (.A1(n_11778_o_0),
    .A2(n_11820_o_0),
    .B(n_11821_o_0),
    .Y(n_11822_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11823 (.A1(n_11818_o_0),
    .A2(n_11819_o_0),
    .B(n_11751_o_0),
    .C(n_11822_o_0),
    .Y(n_11823_o_0));
 OAI211xp5_ASAP7_75t_R n_11824 (.A1(n_11699_o_0),
    .A2(n_11700_o_0),
    .B(n_11752_o_0),
    .C(n_11706_o_0),
    .Y(n_11824_o_0));
 NAND3xp33_ASAP7_75t_R n_11825 (.A(n_11824_o_0),
    .B(n_11773_o_0),
    .C(n_11733_o_0),
    .Y(n_11825_o_0));
 NOR2xp33_ASAP7_75t_R n_11826 (.A(n_11733_o_0),
    .B(n_11707_o_0),
    .Y(n_11826_o_0));
 AOI21xp33_ASAP7_75t_R n_11827 (.A1(n_11778_o_0),
    .A2(n_11826_o_0),
    .B(n_11782_o_0),
    .Y(n_11827_o_0));
 OAI21xp33_ASAP7_75t_R n_11828 (.A1(n_11751_o_0),
    .A2(n_11825_o_0),
    .B(n_11827_o_0),
    .Y(n_11828_o_0));
 NOR2xp33_ASAP7_75t_R n_11829 (.A(n_1858_o_0),
    .B(n_11680_o_0),
    .Y(n_11829_o_0));
 INVx1_ASAP7_75t_R n_1183 (.A(n_1182_o_0),
    .Y(n_1183_o_0));
 INVx1_ASAP7_75t_R n_11830 (.A(n_11681_o_0),
    .Y(n_11830_o_0));
 NOR2xp33_ASAP7_75t_R n_11831 (.A(n_11829_o_0),
    .B(n_11830_o_0),
    .Y(n_11831_o_0));
 AOI31xp33_ASAP7_75t_R n_11832 (.A1(n_11688_o_0),
    .A2(n_11823_o_0),
    .A3(n_11828_o_0),
    .B(n_11831_o_0),
    .Y(n_11832_o_0));
 OAI21xp33_ASAP7_75t_R n_11833 (.A1(n_11799_o_0),
    .A2(n_11815_o_0),
    .B(n_11832_o_0),
    .Y(n_11833_o_0));
 OAI21xp33_ASAP7_75t_R n_11834 (.A1(n_11681_o_1),
    .A2(n_11802_o_0),
    .B(n_11833_o_0),
    .Y(n_11834_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11835 (.A1(n_11671_o_0),
    .A2(net),
    .B(n_11672_o_0),
    .C(_00962_),
    .Y(n_11835_o_0));
 NOR3xp33_ASAP7_75t_R n_11836 (.A(n_11816_o_0),
    .B(n_11751_o_0),
    .C(n_11766_o_0),
    .Y(n_11836_o_0));
 NAND4xp25_ASAP7_75t_R n_11837 (.A(n_11789_o_0),
    .B(n_11766_o_0),
    .C(n_11707_o_0),
    .D(n_11752_o_0),
    .Y(n_11837_o_0));
 AOI21xp33_ASAP7_75t_R n_11838 (.A1(n_11837_o_0),
    .A2(n_11786_o_0),
    .B(n_11761_o_0),
    .Y(n_11838_o_0));
 OAI21xp33_ASAP7_75t_R n_11839 (.A1(n_11836_o_0),
    .A2(n_11838_o_0),
    .B(n_11681_o_1),
    .Y(n_11839_o_0));
 OAI31xp33_ASAP7_75t_R n_1184 (.A1(n_878_o_0),
    .A2(n_907_o_0),
    .A3(n_887_o_0),
    .B(n_1094_o_0),
    .Y(n_1184_o_0));
 NOR2xp33_ASAP7_75t_R n_11840 (.A(n_11766_o_0),
    .B(n_11748_o_0),
    .Y(n_11840_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11841 (.A1(n_11764_o_0),
    .A2(n_11766_o_0),
    .B(n_11840_o_0),
    .C(n_11789_o_0),
    .Y(n_11841_o_0));
 INVx1_ASAP7_75t_R n_11842 (.A(n_11841_o_0),
    .Y(n_11842_o_0));
 NAND2xp33_ASAP7_75t_R n_11843 (.A(n_11752_o_0),
    .B(n_11748_o_0),
    .Y(n_11843_o_0));
 OAI21xp33_ASAP7_75t_R n_11844 (.A1(n_11766_o_0),
    .A2(n_11752_o_0),
    .B(n_11778_o_0),
    .Y(n_11844_o_0));
 INVx2_ASAP7_75t_R n_11845 (.A(n_11782_o_0),
    .Y(n_11845_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11846 (.A1(n_11766_o_0),
    .A2(n_11843_o_0),
    .B(n_11844_o_0),
    .C(n_11845_o_0),
    .Y(n_11846_o_0));
 NOR3xp33_ASAP7_75t_R n_11847 (.A(n_11707_o_0),
    .B(n_11766_o_0),
    .C(n_11752_o_0),
    .Y(n_11847_o_0));
 NOR2xp33_ASAP7_75t_R n_11848 (.A(n_11733_o_0),
    .B(n_11748_o_0),
    .Y(n_11848_o_0));
 NOR3xp33_ASAP7_75t_R n_11849 (.A(n_11847_o_0),
    .B(n_11848_o_0),
    .C(n_11751_o_0),
    .Y(n_11849_o_0));
 AOI21xp33_ASAP7_75t_R n_1185 (.A1(n_891_o_0),
    .A2(n_1184_o_0),
    .B(n_904_o_0),
    .Y(n_1185_o_0));
 OA21x2_ASAP7_75t_R n_11850 (.A1(n_11846_o_0),
    .A2(n_11849_o_0),
    .B(n_11831_o_0),
    .Y(n_11850_o_0));
 OAI21xp33_ASAP7_75t_R n_11851 (.A1(n_11796_o_0),
    .A2(n_11842_o_0),
    .B(n_11850_o_0),
    .Y(n_11851_o_0));
 NOR3xp33_ASAP7_75t_R n_11852 (.A(n_11707_o_0),
    .B(n_11719_o_0),
    .C(n_11733_o_0),
    .Y(n_11852_o_0));
 NOR2xp33_ASAP7_75t_R n_11853 (.A(n_11789_o_0),
    .B(n_11852_o_0),
    .Y(n_11853_o_0));
 NAND2xp33_ASAP7_75t_R n_11854 (.A(n_11733_o_0),
    .B(n_11719_o_0),
    .Y(n_11854_o_0));
 NAND3xp33_ASAP7_75t_R n_11855 (.A(n_11853_o_0),
    .B(n_11854_o_0),
    .C(n_11761_o_0),
    .Y(n_11855_o_0));
 AOI31xp33_ASAP7_75t_R n_11856 (.A1(n_11839_o_0),
    .A2(n_11851_o_0),
    .A3(n_11855_o_0),
    .B(n_11689_o_0),
    .Y(n_11856_o_0));
 INVx1_ASAP7_75t_R n_11857 (.A(n_11831_o_0),
    .Y(n_11857_o_0));
 NOR3xp33_ASAP7_75t_R n_11858 (.A(n_11707_o_0),
    .B(n_11766_o_0),
    .C(n_11752_o_0),
    .Y(n_11858_o_0));
 NOR2xp33_ASAP7_75t_R n_11859 (.A(n_11778_o_0),
    .B(n_11858_o_0),
    .Y(n_11859_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_1186 (.A1(n_878_o_0),
    .A2(n_1180_o_0),
    .B(n_1183_o_0),
    .C(n_1185_o_0),
    .D(n_930_o_0),
    .Y(n_1186_o_0));
 AOI21xp33_ASAP7_75t_R n_11860 (.A1(n_11773_o_0),
    .A2(n_11824_o_0),
    .B(n_11733_o_0),
    .Y(n_11860_o_0));
 AOI21xp33_ASAP7_75t_R n_11861 (.A1(n_11752_o_0),
    .A2(n_11748_o_0),
    .B(n_11766_o_0),
    .Y(n_11861_o_0));
 OAI31xp33_ASAP7_75t_R n_11862 (.A1(n_11789_o_0),
    .A2(n_11860_o_0),
    .A3(n_11861_o_0),
    .B(n_11796_o_0),
    .Y(n_11862_o_0));
 NOR2xp33_ASAP7_75t_R n_11863 (.A(n_11752_o_0),
    .B(n_11707_o_0),
    .Y(n_11863_o_0));
 OAI21xp33_ASAP7_75t_R n_11864 (.A1(n_11733_o_0),
    .A2(n_11863_o_0),
    .B(n_11778_o_0),
    .Y(n_11864_o_0));
 AOI21xp33_ASAP7_75t_R n_11865 (.A1(n_11733_o_0),
    .A2(n_11719_o_0),
    .B(n_11751_o_0),
    .Y(n_11865_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11866 (.A1(_00960_),
    .A2(n_11759_o_0),
    .B(n_11760_o_0),
    .C(n_11865_o_0),
    .Y(n_11866_o_0));
 OAI21xp33_ASAP7_75t_R n_11867 (.A1(n_11847_o_0),
    .A2(n_11864_o_0),
    .B(n_11866_o_0),
    .Y(n_11867_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11868 (.A1(n_11859_o_0),
    .A2(n_11811_o_0),
    .B(n_11862_o_0),
    .C(n_11867_o_0),
    .Y(n_11868_o_0));
 AOI21xp33_ASAP7_75t_R n_11869 (.A1(n_11719_o_0),
    .A2(n_11707_o_0),
    .B(n_11766_o_0),
    .Y(n_11869_o_0));
 OA21x2_ASAP7_75t_R n_1187 (.A1(n_1177_o_0),
    .A2(n_1179_o_0),
    .B(n_1186_o_0),
    .Y(n_1187_o_0));
 INVx1_ASAP7_75t_R n_11870 (.A(n_11869_o_0),
    .Y(n_11870_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11871 (.A1(n_11807_o_0),
    .A2(n_11870_o_0),
    .B(n_11751_o_0),
    .C(n_11864_o_0),
    .Y(n_11871_o_0));
 INVx1_ASAP7_75t_R n_11872 (.A(n_11825_o_0),
    .Y(n_11872_o_0));
 NOR2xp33_ASAP7_75t_R n_11873 (.A(n_11733_o_0),
    .B(n_11707_o_0),
    .Y(n_11873_o_0));
 NAND3xp33_ASAP7_75t_R n_11874 (.A(n_11809_o_0),
    .B(n_11811_o_0),
    .C(n_11751_o_0),
    .Y(n_11874_o_0));
 OAI311xp33_ASAP7_75t_R n_11875 (.A1(n_11778_o_0),
    .A2(n_11872_o_0),
    .A3(n_11873_o_0),
    .B1(n_11874_o_0),
    .C1(n_11782_o_0),
    .Y(n_11875_o_0));
 OAI211xp5_ASAP7_75t_R n_11876 (.A1(n_11782_o_0),
    .A2(n_11871_o_0),
    .B(n_11875_o_0),
    .C(n_11681_o_1),
    .Y(n_11876_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11877 (.A1(n_11857_o_0),
    .A2(n_11868_o_0),
    .B(n_11876_o_0),
    .C(n_11799_o_0),
    .Y(n_11877_o_0));
 AOI211xp5_ASAP7_75t_R n_11878 (.A1(n_11674_o_0),
    .A2(n_11835_o_0),
    .B(n_11856_o_0),
    .C(n_11877_o_0),
    .Y(n_11878_o_0));
 AOI21xp33_ASAP7_75t_R n_11879 (.A1(n_11675_o_0),
    .A2(n_11834_o_0),
    .B(n_11878_o_0),
    .Y(n_11879_o_0));
 AOI21xp33_ASAP7_75t_R n_1188 (.A1(n_930_o_0),
    .A2(n_1175_o_0),
    .B(n_1187_o_0),
    .Y(n_1188_o_0));
 INVx1_ASAP7_75t_R n_11880 (.A(n_11861_o_0),
    .Y(n_11880_o_0));
 NAND2xp33_ASAP7_75t_R n_11881 (.A(n_11766_o_0),
    .B(n_11707_o_0),
    .Y(n_11881_o_0));
 NAND3xp33_ASAP7_75t_R n_11882 (.A(n_11880_o_0),
    .B(n_11881_o_0),
    .C(n_11751_o_0),
    .Y(n_11882_o_0));
 INVx1_ASAP7_75t_R n_11883 (.A(n_11882_o_0),
    .Y(n_11883_o_0));
 OAI21xp33_ASAP7_75t_R n_11884 (.A1(n_11741_o_0),
    .A2(n_11777_o_0),
    .B(n_11766_o_0),
    .Y(n_11884_o_0));
 AOI21xp33_ASAP7_75t_R n_11885 (.A1(net76),
    .A2(n_11752_o_0),
    .B(n_11884_o_0),
    .Y(n_11885_o_0));
 NOR3xp33_ASAP7_75t_R n_11886 (.A(n_11883_o_0),
    .B(n_11799_o_0),
    .C(n_11885_o_0),
    .Y(n_11886_o_0));
 INVx1_ASAP7_75t_R n_11887 (.A(n_11788_o_0),
    .Y(n_11887_o_0));
 NOR3xp33_ASAP7_75t_R n_11888 (.A(n_11707_o_0),
    .B(n_11766_o_0),
    .C(n_11752_o_0),
    .Y(n_11888_o_0));
 AOI211xp5_ASAP7_75t_R n_11889 (.A1(n_11774_o_0),
    .A2(n_11766_o_0),
    .B(n_11888_o_0),
    .C(n_11789_o_0),
    .Y(n_11889_o_0));
 NAND2xp33_ASAP7_75t_R n_1189 (.A(n_877_o_0),
    .B(n_861_o_0),
    .Y(n_1189_o_0));
 AOI31xp33_ASAP7_75t_R n_11890 (.A1(n_11743_o_0),
    .A2(n_11887_o_0),
    .A3(n_11753_o_0),
    .B(n_11889_o_0),
    .Y(n_11890_o_0));
 OAI21xp33_ASAP7_75t_R n_11891 (.A1(n_11798_o_0),
    .A2(n_11890_o_0),
    .B(n_11796_o_0),
    .Y(n_11891_o_0));
 NAND2xp33_ASAP7_75t_R n_11892 (.A(n_11752_o_0),
    .B(n_11748_o_0),
    .Y(n_11892_o_0));
 AOI21xp33_ASAP7_75t_R n_11893 (.A1(n_11733_o_0),
    .A2(n_11774_o_0),
    .B(n_11744_o_0),
    .Y(n_11893_o_0));
 AOI31xp33_ASAP7_75t_R n_11894 (.A1(n_11751_o_0),
    .A2(n_11811_o_0),
    .A3(n_11892_o_0),
    .B(n_11893_o_0),
    .Y(n_11894_o_0));
 NOR2xp33_ASAP7_75t_R n_11895 (.A(n_11733_o_0),
    .B(n_11774_o_0),
    .Y(n_11895_o_0));
 NOR3xp33_ASAP7_75t_R n_11896 (.A(n_11707_o_0),
    .B(n_11719_o_0),
    .C(n_11766_o_0),
    .Y(n_11896_o_0));
 NOR2xp33_ASAP7_75t_R n_11897 (.A(n_11733_o_0),
    .B(n_11751_o_0),
    .Y(n_11897_o_0));
 INVx1_ASAP7_75t_R n_11898 (.A(n_11897_o_0),
    .Y(n_11898_o_0));
 OAI321xp33_ASAP7_75t_R n_11899 (.A1(n_11895_o_0),
    .A2(n_11896_o_0),
    .A3(n_11743_o_0),
    .B1(n_11898_o_0),
    .B2(n_11816_o_0),
    .C(n_11689_o_0),
    .Y(n_11899_o_0));
 NOR2xp33_ASAP7_75t_R n_1190 (.A(n_878_o_0),
    .B(n_956_o_0),
    .Y(n_1190_o_0));
 OAI211xp5_ASAP7_75t_R n_11900 (.A1(n_11894_o_0),
    .A2(n_11798_o_0),
    .B(n_11899_o_0),
    .C(n_11782_o_0),
    .Y(n_11900_o_0));
 OAI21xp33_ASAP7_75t_R n_11901 (.A1(n_11886_o_0),
    .A2(n_11891_o_0),
    .B(n_11900_o_0),
    .Y(n_11901_o_0));
 INVx1_ASAP7_75t_R n_11902 (.A(n_11818_o_0),
    .Y(n_11902_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11903 (.A1(n_11824_o_0),
    .A2(n_11773_o_0),
    .B(n_11766_o_0),
    .C(n_11778_o_0),
    .Y(n_11903_o_0));
 AO21x1_ASAP7_75t_R n_11904 (.A1(n_11766_o_0),
    .A2(n_11843_o_0),
    .B(n_11903_o_0),
    .Y(n_11904_o_0));
 INVx1_ASAP7_75t_R n_11905 (.A(n_11904_o_0),
    .Y(n_11905_o_0));
 NOR2xp33_ASAP7_75t_R n_11906 (.A(n_11766_o_0),
    .B(n_11707_o_0),
    .Y(n_11906_o_0));
 NOR2xp33_ASAP7_75t_R n_11907 (.A(n_11766_o_0),
    .B(n_11751_o_0),
    .Y(n_11907_o_0));
 AOI21xp33_ASAP7_75t_R n_11908 (.A1(n_11863_o_0),
    .A2(n_11907_o_0),
    .B(n_11782_o_0),
    .Y(n_11908_o_0));
 OAI211xp5_ASAP7_75t_R n_11909 (.A1(n_11906_o_0),
    .A2(n_11743_o_0),
    .B(n_11908_o_0),
    .C(n_11881_o_0),
    .Y(n_11909_o_0));
 NOR2xp33_ASAP7_75t_R n_1191 (.A(n_1041_o_0),
    .B(n_1190_o_0),
    .Y(n_1191_o_0));
 OAI31xp33_ASAP7_75t_R n_11910 (.A1(n_11796_o_0),
    .A2(n_11902_o_0),
    .A3(n_11905_o_0),
    .B(n_11909_o_0),
    .Y(n_11910_o_0));
 OAI21xp33_ASAP7_75t_R n_11911 (.A1(n_11689_o_0),
    .A2(n_11910_o_0),
    .B(n_11675_o_0),
    .Y(n_11911_o_0));
 AOI211xp5_ASAP7_75t_R n_11912 (.A1(n_11707_o_0),
    .A2(n_11719_o_0),
    .B(n_11873_o_0),
    .C(n_11778_o_0),
    .Y(n_11912_o_0));
 INVx1_ASAP7_75t_R n_11913 (.A(n_11749_o_0),
    .Y(n_11913_o_0));
 OAI21xp33_ASAP7_75t_R n_11914 (.A1(n_11763_o_0),
    .A2(n_11913_o_0),
    .B(n_11782_o_0),
    .Y(n_11914_o_0));
 NOR2xp33_ASAP7_75t_R n_11915 (.A(n_11752_o_0),
    .B(n_11766_o_0),
    .Y(n_11915_o_0));
 AOI21xp33_ASAP7_75t_R n_11916 (.A1(n_11766_o_0),
    .A2(n_11774_o_0),
    .B(n_11789_o_0),
    .Y(n_11916_o_0));
 INVx1_ASAP7_75t_R n_11917 (.A(n_11916_o_0),
    .Y(n_11917_o_0));
 OAI21xp33_ASAP7_75t_R n_11918 (.A1(n_11733_o_0),
    .A2(n_11863_o_0),
    .B(n_11789_o_0),
    .Y(n_11918_o_0));
 OA21x2_ASAP7_75t_R n_11919 (.A1(n_11918_o_0),
    .A2(n_11820_o_0),
    .B(n_11796_o_0),
    .Y(n_11919_o_0));
 OAI31xp33_ASAP7_75t_R n_1192 (.A1(n_878_o_0),
    .A2(n_907_o_0),
    .A3(n_938_o_0),
    .B(n_891_o_0),
    .Y(n_1192_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11920 (.A1(n_11915_o_0),
    .A2(n_11917_o_0),
    .B(n_11919_o_0),
    .C(n_11688_o_0),
    .Y(n_11920_o_0));
 OA21x2_ASAP7_75t_R n_11921 (.A1(n_11912_o_0),
    .A2(n_11914_o_0),
    .B(n_11920_o_0),
    .Y(n_11921_o_0));
 OAI22xp33_ASAP7_75t_R n_11922 (.A1(n_11901_o_0),
    .A2(n_11675_o_0),
    .B1(n_11911_o_0),
    .B2(n_11921_o_0),
    .Y(n_11922_o_0));
 NAND2xp33_ASAP7_75t_R n_11923 (.A(n_11733_o_0),
    .B(n_11707_o_0),
    .Y(n_11923_o_0));
 INVx1_ASAP7_75t_R n_11924 (.A(n_11864_o_0),
    .Y(n_11924_o_0));
 OAI21xp33_ASAP7_75t_R n_11925 (.A1(n_11792_o_0),
    .A2(n_11744_o_0),
    .B(n_11688_o_0),
    .Y(n_11925_o_0));
 AOI21xp33_ASAP7_75t_R n_11926 (.A1(n_11923_o_0),
    .A2(n_11924_o_0),
    .B(n_11925_o_0),
    .Y(n_11926_o_0));
 INVx1_ASAP7_75t_R n_11927 (.A(n_11858_o_0),
    .Y(n_11927_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11928 (.A1(n_11707_o_0),
    .A2(n_11766_o_0),
    .B(n_11719_o_0),
    .C(n_11778_o_0),
    .Y(n_11928_o_0));
 AOI211xp5_ASAP7_75t_R n_11929 (.A1(n_11853_o_0),
    .A2(n_11927_o_0),
    .B(n_11799_o_0),
    .C(n_11928_o_0),
    .Y(n_11929_o_0));
 AOI21xp33_ASAP7_75t_R n_1193 (.A1(n_878_o_0),
    .A2(net32),
    .B(n_1192_o_0),
    .Y(n_1193_o_0));
 NAND2xp33_ASAP7_75t_R n_11930 (.A(n_11719_o_0),
    .B(n_11707_o_0),
    .Y(n_11930_o_0));
 OAI21xp33_ASAP7_75t_R n_11931 (.A1(n_11719_o_0),
    .A2(n_11766_o_0),
    .B(n_11789_o_0),
    .Y(n_11931_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11932 (.A1(n_11785_o_0),
    .A2(n_11733_o_0),
    .B(n_11743_o_0),
    .C(n_11931_o_0),
    .Y(n_11932_o_0));
 NAND3xp33_ASAP7_75t_R n_11933 (.A(n_11930_o_0),
    .B(n_11751_o_0),
    .C(n_11766_o_0),
    .Y(n_11933_o_0));
 OAI211xp5_ASAP7_75t_R n_11934 (.A1(n_11930_o_0),
    .A2(n_11884_o_0),
    .B(n_11932_o_0),
    .C(n_11933_o_0),
    .Y(n_11934_o_0));
 AOI21xp33_ASAP7_75t_R n_11935 (.A1(n_11766_o_0),
    .A2(n_11843_o_0),
    .B(n_11751_o_0),
    .Y(n_11935_o_0));
 OAI21xp33_ASAP7_75t_R n_11936 (.A1(n_11766_o_0),
    .A2(n_11764_o_0),
    .B(n_11935_o_0),
    .Y(n_11936_o_0));
 OAI311xp33_ASAP7_75t_R n_11937 (.A1(n_11743_o_0),
    .A2(n_11895_o_0),
    .A3(n_11896_o_0),
    .B1(n_11799_o_0),
    .C1(n_11936_o_0),
    .Y(n_11937_o_0));
 OAI211xp5_ASAP7_75t_R n_11938 (.A1(n_11934_o_0),
    .A2(n_11799_o_0),
    .B(n_11937_o_0),
    .C(n_11674_o_1),
    .Y(n_11938_o_0));
 OAI31xp33_ASAP7_75t_R n_11939 (.A1(n_11674_o_1),
    .A2(n_11926_o_0),
    .A3(n_11929_o_0),
    .B(n_11938_o_0),
    .Y(n_11939_o_0));
 AOI311xp33_ASAP7_75t_R n_1194 (.A1(n_1189_o_0),
    .A2(n_1191_o_0),
    .A3(net16),
    .B(n_904_o_0),
    .C(n_1193_o_0),
    .Y(n_1194_o_0));
 NAND2xp33_ASAP7_75t_R n_11940 (.A(n_11733_o_0),
    .B(n_11707_o_0),
    .Y(n_11940_o_0));
 INVx1_ASAP7_75t_R n_11941 (.A(n_11852_o_0),
    .Y(n_11941_o_0));
 NAND3xp33_ASAP7_75t_R n_11942 (.A(n_11941_o_0),
    .B(n_11809_o_0),
    .C(n_11743_o_0),
    .Y(n_11942_o_0));
 INVx1_ASAP7_75t_R n_11943 (.A(n_11942_o_0),
    .Y(n_11943_o_0));
 AOI31xp33_ASAP7_75t_R n_11944 (.A1(n_11751_o_0),
    .A2(n_11799_o_0),
    .A3(n_11940_o_0),
    .B(n_11943_o_0),
    .Y(n_11944_o_0));
 AOI21xp33_ASAP7_75t_R n_11945 (.A1(n_11923_o_0),
    .A2(n_11924_o_0),
    .B(n_11688_o_0),
    .Y(n_11945_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11946 (.A1(n_11733_o_0),
    .A2(n_11764_o_0),
    .B(n_11744_o_0),
    .C(n_11945_o_0),
    .Y(n_11946_o_0));
 OAI31xp33_ASAP7_75t_R n_11947 (.A1(n_11778_o_0),
    .A2(n_11852_o_0),
    .A3(n_11915_o_0),
    .B(n_11688_o_0),
    .Y(n_11947_o_0));
 NAND2xp33_ASAP7_75t_R n_11948 (.A(n_11835_o_0),
    .B(n_11674_o_0),
    .Y(n_11948_o_0));
 OA21x2_ASAP7_75t_R n_11949 (.A1(n_11947_o_0),
    .A2(n_11916_o_0),
    .B(n_11948_o_0),
    .Y(n_11949_o_0));
 NAND3xp33_ASAP7_75t_R n_1195 (.A(n_941_o_0),
    .B(n_990_o_0),
    .C(n_877_o_0),
    .Y(n_1195_o_0));
 AOI21xp33_ASAP7_75t_R n_11950 (.A1(n_11946_o_0),
    .A2(n_11949_o_0),
    .B(n_11845_o_0),
    .Y(n_11950_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11951 (.A1(n_11674_o_1),
    .A2(n_11944_o_0),
    .B(n_11950_o_0),
    .C(n_11681_o_1),
    .Y(n_11951_o_0));
 OAI21xp33_ASAP7_75t_R n_11952 (.A1(n_11761_o_0),
    .A2(n_11939_o_0),
    .B(n_11951_o_0),
    .Y(n_11952_o_0));
 OAI21xp33_ASAP7_75t_R n_11953 (.A1(n_11831_o_0),
    .A2(n_11922_o_0),
    .B(n_11952_o_0),
    .Y(n_11953_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11954 (.A1(n_11733_o_0),
    .A2(n_11816_o_0),
    .B(n_11806_o_0),
    .C(n_11751_o_0),
    .Y(n_11954_o_0));
 OAI31xp33_ASAP7_75t_R n_11955 (.A1(n_11778_o_0),
    .A2(n_11872_o_0),
    .A3(n_11873_o_0),
    .B(n_11954_o_0),
    .Y(n_11955_o_0));
 NOR2xp33_ASAP7_75t_R n_11956 (.A(n_11733_o_0),
    .B(n_11707_o_0),
    .Y(n_11956_o_0));
 NOR3xp33_ASAP7_75t_R n_11957 (.A(n_11847_o_0),
    .B(n_11743_o_0),
    .C(n_11956_o_0),
    .Y(n_11957_o_0));
 OAI21xp33_ASAP7_75t_R n_11958 (.A1(n_11861_o_0),
    .A2(n_11918_o_0),
    .B(n_11688_o_0),
    .Y(n_11958_o_0));
 NAND2xp33_ASAP7_75t_R n_11959 (.A(n_11761_o_0),
    .B(n_11799_o_0),
    .Y(n_11959_o_0));
 AOI211xp5_ASAP7_75t_R n_1196 (.A1(n_916_o_0),
    .A2(n_877_o_0),
    .B(net14),
    .C(n_1012_o_0),
    .Y(n_1196_o_0));
 OAI21xp33_ASAP7_75t_R n_11960 (.A1(n_11957_o_0),
    .A2(n_11958_o_0),
    .B(n_11959_o_0),
    .Y(n_11960_o_0));
 NAND2xp33_ASAP7_75t_R n_11961 (.A(n_11752_o_0),
    .B(n_11766_o_0),
    .Y(n_11961_o_0));
 AOI311xp33_ASAP7_75t_R n_11962 (.A1(n_11766_o_0),
    .A2(n_11824_o_0),
    .A3(n_11773_o_0),
    .B(n_11778_o_0),
    .C(n_11840_o_0),
    .Y(n_11962_o_0));
 AOI31xp33_ASAP7_75t_R n_11963 (.A1(n_11961_o_0),
    .A2(n_11751_o_0),
    .A3(n_11819_o_0),
    .B(n_11962_o_0),
    .Y(n_11963_o_0));
 AO21x1_ASAP7_75t_R n_11964 (.A1(n_11843_o_0),
    .A2(n_11766_o_0),
    .B(n_11896_o_0),
    .Y(n_11964_o_0));
 NAND2xp33_ASAP7_75t_R n_11965 (.A(n_11761_o_0),
    .B(n_11689_o_0),
    .Y(n_11965_o_0));
 INVx1_ASAP7_75t_R n_11966 (.A(n_11965_o_0),
    .Y(n_11966_o_0));
 OAI221xp5_ASAP7_75t_R n_11967 (.A1(n_11743_o_0),
    .A2(n_11964_o_0),
    .B1(n_11751_o_0),
    .B2(n_11847_o_0),
    .C(n_11966_o_0),
    .Y(n_11967_o_0));
 OAI31xp33_ASAP7_75t_R n_11968 (.A1(n_11688_o_0),
    .A2(n_11782_o_0),
    .A3(n_11963_o_0),
    .B(n_11967_o_0),
    .Y(n_11968_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11969 (.A1(n_11845_o_0),
    .A2(n_11955_o_0),
    .B(n_11960_o_0),
    .C(n_11968_o_0),
    .Y(n_11969_o_0));
 AOI311xp33_ASAP7_75t_R n_1197 (.A1(net15),
    .A2(n_959_o_0),
    .A3(n_1195_o_0),
    .B(n_903_o_0),
    .C(n_1196_o_0),
    .Y(n_1197_o_0));
 OAI31xp33_ASAP7_75t_R n_11970 (.A1(n_11707_o_0),
    .A2(n_11766_o_0),
    .A3(n_11751_o_0),
    .B(n_11845_o_0),
    .Y(n_11970_o_0));
 OAI22xp33_ASAP7_75t_R n_11971 (.A1(n_11858_o_0),
    .A2(n_11778_o_0),
    .B1(n_11789_o_0),
    .B2(n_11826_o_0),
    .Y(n_11971_o_0));
 OAI22xp33_ASAP7_75t_R n_11972 (.A1(n_11957_o_0),
    .A2(n_11970_o_0),
    .B1(n_11971_o_0),
    .B2(n_11845_o_0),
    .Y(n_11972_o_0));
 OAI21xp33_ASAP7_75t_R n_11973 (.A1(n_11733_o_0),
    .A2(n_11719_o_0),
    .B(n_11751_o_0),
    .Y(n_11973_o_0));
 OA21x2_ASAP7_75t_R n_11974 (.A1(n_11973_o_0),
    .A2(n_11765_o_0),
    .B(n_11796_o_0),
    .Y(n_11974_o_0));
 OAI21xp33_ASAP7_75t_R n_11975 (.A1(n_11852_o_0),
    .A2(n_11810_o_0),
    .B(n_11974_o_0),
    .Y(n_11975_o_0));
 AOI21xp33_ASAP7_75t_R n_11976 (.A1(n_11930_o_0),
    .A2(n_11897_o_0),
    .B(n_11796_o_0),
    .Y(n_11976_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_11977 (.A1(n_11733_o_0),
    .A2(n_11816_o_0),
    .B(n_11786_o_0),
    .C(n_11976_o_0),
    .Y(n_11977_o_0));
 AOI31xp33_ASAP7_75t_R n_11978 (.A1(n_11798_o_0),
    .A2(n_11975_o_0),
    .A3(n_11977_o_0),
    .B(n_11831_o_0),
    .Y(n_11978_o_0));
 OAI21xp33_ASAP7_75t_R n_11979 (.A1(n_11689_o_0),
    .A2(n_11972_o_0),
    .B(n_11978_o_0),
    .Y(n_11979_o_0));
 NAND2xp33_ASAP7_75t_R n_1198 (.A(n_1182_o_0),
    .B(n_1153_o_0),
    .Y(n_1198_o_0));
 OAI21xp33_ASAP7_75t_R n_11980 (.A1(n_11681_o_1),
    .A2(n_11969_o_0),
    .B(n_11979_o_0),
    .Y(n_11980_o_0));
 INVx1_ASAP7_75t_R n_11981 (.A(n_11744_o_0),
    .Y(n_11981_o_0));
 OAI21xp33_ASAP7_75t_R n_11982 (.A1(n_11766_o_0),
    .A2(n_11767_o_0),
    .B(n_11981_o_0),
    .Y(n_11982_o_0));
 OAI211xp5_ASAP7_75t_R n_11983 (.A1(n_11895_o_0),
    .A2(n_11903_o_0),
    .B(n_11982_o_0),
    .C(n_11782_o_0),
    .Y(n_11983_o_0));
 OAI21xp33_ASAP7_75t_R n_11984 (.A1(net76),
    .A2(n_11766_o_0),
    .B(n_11751_o_0),
    .Y(n_11984_o_0));
 NOR2xp33_ASAP7_75t_R n_11985 (.A(n_11733_o_0),
    .B(n_11767_o_0),
    .Y(n_11985_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_11986 (.A1(n_11766_o_0),
    .A2(n_11843_o_0),
    .B(n_11981_o_0),
    .C(n_11761_o_0),
    .Y(n_11986_o_0));
 OAI21xp33_ASAP7_75t_R n_11987 (.A1(n_11984_o_0),
    .A2(n_11985_o_0),
    .B(n_11986_o_0),
    .Y(n_11987_o_0));
 NOR2xp33_ASAP7_75t_R n_11988 (.A(n_11766_o_0),
    .B(n_11843_o_0),
    .Y(n_11988_o_0));
 NOR2xp33_ASAP7_75t_R n_11989 (.A(n_11985_o_0),
    .B(n_11988_o_0),
    .Y(n_11989_o_0));
 OAI31xp33_ASAP7_75t_R n_1199 (.A1(net16),
    .A2(n_911_o_0),
    .A3(n_976_o_0),
    .B(n_1198_o_0),
    .Y(n_1199_o_0));
 AOI211xp5_ASAP7_75t_R n_11990 (.A1(n_11766_o_0),
    .A2(n_11752_o_0),
    .B(n_11888_o_0),
    .C(n_11789_o_0),
    .Y(n_11990_o_0));
 AOI21xp33_ASAP7_75t_R n_11991 (.A1(n_11743_o_0),
    .A2(n_11989_o_0),
    .B(n_11990_o_0),
    .Y(n_11991_o_0));
 AOI22xp33_ASAP7_75t_R n_11992 (.A1(n_11897_o_0),
    .A2(n_11803_o_0),
    .B1(n_11907_o_0),
    .B2(n_11863_o_0),
    .Y(n_11992_o_0));
 OAI211xp5_ASAP7_75t_R n_11993 (.A1(n_11719_o_0),
    .A2(n_11766_o_0),
    .B(n_11778_o_0),
    .C(net76),
    .Y(n_11993_o_0));
 NOR2xp33_ASAP7_75t_R n_11994 (.A(n_11782_o_0),
    .B(n_11798_o_0),
    .Y(n_11994_o_0));
 AOI31xp33_ASAP7_75t_R n_11995 (.A1(n_11799_o_0),
    .A2(n_11992_o_0),
    .A3(n_11993_o_0),
    .B(n_11994_o_0),
    .Y(n_11995_o_0));
 AOI21xp33_ASAP7_75t_R n_11996 (.A1(n_11796_o_0),
    .A2(n_11991_o_0),
    .B(n_11995_o_0),
    .Y(n_11996_o_0));
 AOI31xp33_ASAP7_75t_R n_11997 (.A1(n_11689_o_0),
    .A2(n_11983_o_0),
    .A3(n_11987_o_0),
    .B(n_11996_o_0),
    .Y(n_11997_o_0));
 INVx1_ASAP7_75t_R n_11998 (.A(n_11873_o_0),
    .Y(n_11998_o_0));
 AOI21xp33_ASAP7_75t_R n_11999 (.A1(n_11707_o_0),
    .A2(n_11719_o_0),
    .B(n_11789_o_0),
    .Y(n_11999_o_0));
 NAND3xp33_ASAP7_75t_R n_1200 (.A(n_953_o_0),
    .B(n_1005_o_0),
    .C(n_878_o_0),
    .Y(n_1200_o_0));
 AOI21xp33_ASAP7_75t_R n_12000 (.A1(n_11998_o_0),
    .A2(n_11999_o_0),
    .B(n_11845_o_0),
    .Y(n_12000_o_0));
 INVx1_ASAP7_75t_R n_12001 (.A(n_12000_o_0),
    .Y(n_12001_o_0));
 AOI21xp33_ASAP7_75t_R n_12002 (.A1(n_11752_o_0),
    .A2(n_11707_o_0),
    .B(n_11733_o_0),
    .Y(n_12002_o_0));
 NOR2xp33_ASAP7_75t_R n_12003 (.A(n_11778_o_0),
    .B(n_11873_o_0),
    .Y(n_12003_o_0));
 OAI21xp33_ASAP7_75t_R n_12004 (.A1(n_11766_o_0),
    .A2(n_11764_o_0),
    .B(n_12003_o_0),
    .Y(n_12004_o_0));
 OAI31xp33_ASAP7_75t_R n_12005 (.A1(n_11789_o_0),
    .A2(n_11872_o_0),
    .A3(n_12002_o_0),
    .B(n_12004_o_0),
    .Y(n_12005_o_0));
 AOI21xp33_ASAP7_75t_R n_12006 (.A1(n_11845_o_0),
    .A2(n_12005_o_0),
    .B(n_11689_o_0),
    .Y(n_12006_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12007 (.A1(n_11743_o_0),
    .A2(n_11940_o_0),
    .B(n_12001_o_0),
    .C(n_12006_o_0),
    .Y(n_12007_o_0));
 AOI211xp5_ASAP7_75t_R n_12008 (.A1(n_11785_o_0),
    .A2(n_11733_o_0),
    .B(n_11751_o_0),
    .C(n_11956_o_0),
    .Y(n_12008_o_0));
 NAND3xp33_ASAP7_75t_R n_12009 (.A(n_11923_o_0),
    .B(n_11805_o_0),
    .C(n_11778_o_0),
    .Y(n_12009_o_0));
 NOR2xp33_ASAP7_75t_R n_1201 (.A(n_913_o_0),
    .B(n_878_o_0),
    .Y(n_1201_o_0));
 INVx1_ASAP7_75t_R n_12010 (.A(n_12009_o_0),
    .Y(n_12010_o_0));
 OAI321xp33_ASAP7_75t_R n_12011 (.A1(n_11707_o_0),
    .A2(n_11751_o_0),
    .A3(n_11733_o_0),
    .B1(n_11806_o_0),
    .B2(n_11903_o_0),
    .C(n_11761_o_0),
    .Y(n_12011_o_0));
 OAI31xp33_ASAP7_75t_R n_12012 (.A1(n_11782_o_0),
    .A2(n_12008_o_0),
    .A3(n_12010_o_0),
    .B(n_12011_o_0),
    .Y(n_12012_o_0));
 OA21x2_ASAP7_75t_R n_12013 (.A1(n_12012_o_0),
    .A2(n_11799_o_0),
    .B(n_11857_o_0),
    .Y(n_12013_o_0));
 AOI21xp33_ASAP7_75t_R n_12014 (.A1(n_12007_o_0),
    .A2(n_12013_o_0),
    .B(n_11675_o_0),
    .Y(n_12014_o_0));
 OAI21xp33_ASAP7_75t_R n_12015 (.A1(n_11681_o_1),
    .A2(n_11997_o_0),
    .B(n_12014_o_0),
    .Y(n_12015_o_0));
 OAI21xp33_ASAP7_75t_R n_12016 (.A1(n_11948_o_0),
    .A2(n_11980_o_0),
    .B(n_12015_o_0),
    .Y(n_12016_o_0));
 OAI311xp33_ASAP7_75t_R n_12017 (.A1(n_11778_o_0),
    .A2(n_11860_o_0),
    .A3(n_11787_o_0),
    .B1(n_11796_o_0),
    .C1(n_11754_o_0),
    .Y(n_12017_o_0));
 NAND3xp33_ASAP7_75t_R n_12018 (.A(n_11767_o_0),
    .B(n_11751_o_0),
    .C(n_11766_o_0),
    .Y(n_12018_o_0));
 NAND4xp25_ASAP7_75t_R n_12019 (.A(n_11743_o_0),
    .B(n_11824_o_0),
    .C(n_11773_o_0),
    .D(n_11733_o_0),
    .Y(n_12019_o_0));
 AOI211xp5_ASAP7_75t_R n_1202 (.A1(n_990_o_0),
    .A2(n_878_o_0),
    .B(n_1201_o_0),
    .C(n_829_o_0),
    .Y(n_1202_o_0));
 OAI211xp5_ASAP7_75t_R n_12020 (.A1(n_11913_o_0),
    .A2(n_11763_o_0),
    .B(n_12018_o_0),
    .C(n_12019_o_0),
    .Y(n_12020_o_0));
 OAI21xp33_ASAP7_75t_R n_12021 (.A1(n_11885_o_0),
    .A2(n_12020_o_0),
    .B(n_11761_o_0),
    .Y(n_12021_o_0));
 AOI21xp33_ASAP7_75t_R n_12022 (.A1(n_12017_o_0),
    .A2(n_12021_o_0),
    .B(n_11688_o_0),
    .Y(n_12022_o_0));
 INVx1_ASAP7_75t_R n_12023 (.A(n_11787_o_0),
    .Y(n_12023_o_0));
 AOI21xp33_ASAP7_75t_R n_12024 (.A1(n_12023_o_0),
    .A2(n_11795_o_0),
    .B(n_11761_o_0),
    .Y(n_12024_o_0));
 OAI21xp33_ASAP7_75t_R n_12025 (.A1(n_11744_o_0),
    .A2(n_11913_o_0),
    .B(n_11782_o_0),
    .Y(n_12025_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12026 (.A1(n_11751_o_0),
    .A2(n_11927_o_0),
    .B(n_12025_o_0),
    .C(n_11799_o_0),
    .Y(n_12026_o_0));
 AOI21xp33_ASAP7_75t_R n_12027 (.A1(n_12024_o_0),
    .A2(n_11882_o_0),
    .B(n_12026_o_0),
    .Y(n_12027_o_0));
 NOR3xp33_ASAP7_75t_R n_12028 (.A(n_12022_o_0),
    .B(n_12027_o_0),
    .C(n_11675_o_0),
    .Y(n_12028_o_0));
 AOI21xp33_ASAP7_75t_R n_12029 (.A1(n_11766_o_0),
    .A2(n_11930_o_0),
    .B(n_11903_o_0),
    .Y(n_12029_o_0));
 AOI31xp33_ASAP7_75t_R n_1203 (.A1(n_1002_o_0),
    .A2(n_1200_o_0),
    .A3(net16),
    .B(n_1202_o_0),
    .Y(n_1203_o_0));
 AOI21xp33_ASAP7_75t_R n_12030 (.A1(n_11766_o_0),
    .A2(n_11767_o_0),
    .B(n_11931_o_0),
    .Y(n_12030_o_0));
 NAND2xp33_ASAP7_75t_R n_12031 (.A(n_11766_o_0),
    .B(n_11843_o_0),
    .Y(n_12031_o_0));
 AOI21xp33_ASAP7_75t_R n_12032 (.A1(n_11733_o_0),
    .A2(n_11816_o_0),
    .B(n_11743_o_0),
    .Y(n_12032_o_0));
 AO21x1_ASAP7_75t_R n_12033 (.A1(n_12031_o_0),
    .A2(n_12032_o_0),
    .B(n_11845_o_0),
    .Y(n_12033_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12034 (.A1(n_11766_o_0),
    .A2(net76),
    .B(n_11795_o_0),
    .C(n_12033_o_0),
    .Y(n_12034_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12035 (.A1(n_12029_o_0),
    .A2(n_12030_o_0),
    .B(n_11796_o_0),
    .C(n_12034_o_0),
    .Y(n_12035_o_0));
 INVx1_ASAP7_75t_R n_12036 (.A(n_11763_o_0),
    .Y(n_12036_o_0));
 AO21x1_ASAP7_75t_R n_12037 (.A1(n_11774_o_0),
    .A2(n_12036_o_0),
    .B(n_11925_o_0),
    .Y(n_12037_o_0));
 OAI21xp33_ASAP7_75t_R n_12038 (.A1(n_11860_o_0),
    .A2(n_11984_o_0),
    .B(n_11782_o_0),
    .Y(n_12038_o_0));
 AOI21xp33_ASAP7_75t_R n_12039 (.A1(n_11981_o_0),
    .A2(n_11749_o_0),
    .B(n_12038_o_0),
    .Y(n_12039_o_0));
 AOI21xp33_ASAP7_75t_R n_1204 (.A1(n_904_o_0),
    .A2(n_1203_o_0),
    .B(n_931_o_0),
    .Y(n_1204_o_0));
 AOI21xp33_ASAP7_75t_R n_12040 (.A1(n_11959_o_0),
    .A2(n_12037_o_0),
    .B(n_12039_o_0),
    .Y(n_12040_o_0));
 AOI211xp5_ASAP7_75t_R n_12041 (.A1(n_12035_o_0),
    .A2(n_11689_o_0),
    .B(n_11948_o_0),
    .C(n_12040_o_0),
    .Y(n_12041_o_0));
 OAI21xp33_ASAP7_75t_R n_12042 (.A1(n_11744_o_0),
    .A2(n_11988_o_0),
    .B(n_11796_o_0),
    .Y(n_12042_o_0));
 INVx1_ASAP7_75t_R n_12043 (.A(n_11959_o_0),
    .Y(n_12043_o_0));
 NOR2xp33_ASAP7_75t_R n_12044 (.A(n_11733_o_0),
    .B(n_11719_o_0),
    .Y(n_12044_o_0));
 OAI31xp33_ASAP7_75t_R n_12045 (.A1(n_11789_o_0),
    .A2(n_11787_o_0),
    .A3(n_12044_o_0),
    .B(n_11942_o_0),
    .Y(n_12045_o_0));
 AOI21xp33_ASAP7_75t_R n_12046 (.A1(n_12043_o_0),
    .A2(n_12045_o_0),
    .B(n_11675_o_0),
    .Y(n_12046_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12047 (.A1(n_11798_o_0),
    .A2(n_12042_o_0),
    .B(n_12046_o_0),
    .C(n_11681_o_1),
    .Y(n_12047_o_0));
 INVx1_ASAP7_75t_R n_12048 (.A(n_11822_o_0),
    .Y(n_12048_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12049 (.A1(n_11733_o_0),
    .A2(n_11767_o_0),
    .B(n_11854_o_0),
    .C(n_11743_o_0),
    .Y(n_12049_o_0));
 OAI21xp33_ASAP7_75t_R n_1205 (.A1(n_904_o_0),
    .A2(n_1199_o_0),
    .B(n_1204_o_0),
    .Y(n_1205_o_0));
 AOI21xp33_ASAP7_75t_R n_12050 (.A1(n_11880_o_0),
    .A2(n_11779_o_0),
    .B(n_12049_o_0),
    .Y(n_12050_o_0));
 AOI21xp33_ASAP7_75t_R n_12051 (.A1(n_11796_o_0),
    .A2(n_12050_o_0),
    .B(n_11688_o_0),
    .Y(n_12051_o_0));
 OAI21xp33_ASAP7_75t_R n_12052 (.A1(n_11912_o_0),
    .A2(n_12048_o_0),
    .B(n_12051_o_0),
    .Y(n_12052_o_0));
 NOR2xp33_ASAP7_75t_R n_12053 (.A(n_11681_o_1),
    .B(n_12052_o_0),
    .Y(n_12053_o_0));
 NAND3xp33_ASAP7_75t_R n_12054 (.A(n_11998_o_0),
    .B(n_11809_o_0),
    .C(n_11743_o_0),
    .Y(n_12054_o_0));
 OAI31xp33_ASAP7_75t_R n_12055 (.A1(n_11743_o_0),
    .A2(n_11785_o_0),
    .A3(n_11763_o_0),
    .B(n_12054_o_0),
    .Y(n_12055_o_0));
 AOI21xp33_ASAP7_75t_R n_12056 (.A1(n_11789_o_0),
    .A2(n_11860_o_0),
    .B(n_11782_o_0),
    .Y(n_12056_o_0));
 OAI22xp33_ASAP7_75t_R n_12057 (.A1(n_12056_o_0),
    .A2(n_11994_o_0),
    .B1(n_11807_o_0),
    .B2(n_11743_o_0),
    .Y(n_12057_o_0));
 AOI21xp33_ASAP7_75t_R n_12058 (.A1(n_11799_o_0),
    .A2(n_12055_o_0),
    .B(n_12057_o_0),
    .Y(n_12058_o_0));
 NAND2xp33_ASAP7_75t_R n_12059 (.A(n_11854_o_0),
    .B(n_11779_o_0),
    .Y(n_12059_o_0));
 OAI311xp33_ASAP7_75t_R n_1206 (.A1(n_930_o_0),
    .A2(n_1194_o_0),
    .A3(n_1197_o_0),
    .B1(n_971_o_0),
    .C1(n_1205_o_0),
    .Y(n_1206_o_0));
 OAI21xp33_ASAP7_75t_R n_12060 (.A1(n_11861_o_0),
    .A2(n_11973_o_0),
    .B(n_12059_o_0),
    .Y(n_12060_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12061 (.A1(n_11733_o_0),
    .A2(n_11767_o_0),
    .B(n_11778_o_0),
    .C(n_11688_o_0),
    .Y(n_12061_o_0));
 AO21x1_ASAP7_75t_R n_12062 (.A1(n_11982_o_0),
    .A2(n_12061_o_0),
    .B(n_11845_o_0),
    .Y(n_12062_o_0));
 AOI21xp33_ASAP7_75t_R n_12063 (.A1(n_11799_o_0),
    .A2(n_12060_o_0),
    .B(n_12062_o_0),
    .Y(n_12063_o_0));
 INVx1_ASAP7_75t_R n_12064 (.A(n_11948_o_0),
    .Y(n_12064_o_0));
 OAI21xp33_ASAP7_75t_R n_12065 (.A1(n_12058_o_0),
    .A2(n_12063_o_0),
    .B(n_12064_o_0),
    .Y(n_12065_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12066 (.A1(n_12047_o_0),
    .A2(n_12052_o_0),
    .B(n_12053_o_0),
    .C(n_12065_o_0),
    .Y(n_12066_o_0));
 OAI31xp33_ASAP7_75t_R n_12067 (.A1(n_11831_o_0),
    .A2(n_12028_o_0),
    .A3(n_12041_o_0),
    .B(n_12066_o_0),
    .Y(n_12067_o_0));
 AOI21xp33_ASAP7_75t_R n_12068 (.A1(n_11778_o_0),
    .A2(n_11792_o_0),
    .B(n_11798_o_0),
    .Y(n_12068_o_0));
 OAI311xp33_ASAP7_75t_R n_12069 (.A1(n_11743_o_0),
    .A2(n_11733_o_0),
    .A3(n_11764_o_0),
    .B1(n_12068_o_0),
    .C1(n_11818_o_0),
    .Y(n_12069_o_0));
 OAI21xp33_ASAP7_75t_R n_1207 (.A1(n_971_o_0),
    .A2(n_1188_o_0),
    .B(n_1206_o_0),
    .Y(n_1207_o_0));
 NOR2xp33_ASAP7_75t_R n_12070 (.A(n_11766_o_0),
    .B(n_11803_o_0),
    .Y(n_12070_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12071 (.A1(n_11766_o_0),
    .A2(n_11785_o_0),
    .B(n_11935_o_0),
    .C(n_11688_o_0),
    .Y(n_12071_o_0));
 OAI31xp33_ASAP7_75t_R n_12072 (.A1(n_11789_o_0),
    .A2(n_12070_o_0),
    .A3(n_11812_o_0),
    .B(n_12071_o_0),
    .Y(n_12072_o_0));
 AND3x1_ASAP7_75t_R n_12073 (.A(n_12069_o_0),
    .B(n_12072_o_0),
    .C(n_11782_o_0),
    .Y(n_12073_o_0));
 NOR3xp33_ASAP7_75t_R n_12074 (.A(n_11774_o_0),
    .B(n_11766_o_0),
    .C(n_11743_o_0),
    .Y(n_12074_o_0));
 NOR3xp33_ASAP7_75t_R n_12075 (.A(n_11836_o_0),
    .B(n_12074_o_0),
    .C(n_11985_o_0),
    .Y(n_12075_o_0));
 INVx1_ASAP7_75t_R n_12076 (.A(n_11812_o_0),
    .Y(n_12076_o_0));
 AOI31xp33_ASAP7_75t_R n_12077 (.A1(n_11751_o_0),
    .A2(n_12076_o_0),
    .A3(n_11923_o_0),
    .B(n_11958_o_0),
    .Y(n_12077_o_0));
 AOI211xp5_ASAP7_75t_R n_12078 (.A1(n_11689_o_0),
    .A2(n_12075_o_0),
    .B(n_12077_o_0),
    .C(n_11761_o_0),
    .Y(n_12078_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12079 (.A1(n_11707_o_0),
    .A2(n_11766_o_0),
    .B(n_11719_o_0),
    .C(n_11751_o_0),
    .Y(n_12079_o_0));
 OAI21xp33_ASAP7_75t_R n_1208 (.A1(n_942_o_0),
    .A2(n_1050_o_0),
    .B(n_904_o_0),
    .Y(n_1208_o_0));
 AOI211xp5_ASAP7_75t_R n_12080 (.A1(n_11719_o_0),
    .A2(n_11766_o_0),
    .B(n_11906_o_0),
    .C(n_11743_o_0),
    .Y(n_12080_o_0));
 AO21x1_ASAP7_75t_R n_12081 (.A1(n_11998_o_0),
    .A2(n_11999_o_0),
    .B(n_11925_o_0),
    .Y(n_12081_o_0));
 OAI31xp33_ASAP7_75t_R n_12082 (.A1(n_11688_o_0),
    .A2(n_12079_o_0),
    .A3(n_12080_o_0),
    .B(n_12081_o_0),
    .Y(n_12082_o_0));
 AOI21xp33_ASAP7_75t_R n_12083 (.A1(n_11870_o_0),
    .A2(n_11998_o_0),
    .B(n_11743_o_0),
    .Y(n_12083_o_0));
 NAND3xp33_ASAP7_75t_R n_12084 (.A(n_11892_o_0),
    .B(n_11881_o_0),
    .C(n_11743_o_0),
    .Y(n_12084_o_0));
 INVx1_ASAP7_75t_R n_12085 (.A(n_12084_o_0),
    .Y(n_12085_o_0));
 NAND3xp33_ASAP7_75t_R n_12086 (.A(n_11804_o_0),
    .B(n_11807_o_0),
    .C(n_11689_o_0),
    .Y(n_12086_o_0));
 OAI31xp33_ASAP7_75t_R n_12087 (.A1(n_11798_o_0),
    .A2(n_12083_o_0),
    .A3(n_12085_o_0),
    .B(n_12086_o_0),
    .Y(n_12087_o_0));
 OAI221xp5_ASAP7_75t_R n_12088 (.A1(n_11845_o_0),
    .A2(n_12082_o_0),
    .B1(n_11761_o_0),
    .B2(n_12087_o_0),
    .C(n_11948_o_0),
    .Y(n_12088_o_0));
 OAI31xp33_ASAP7_75t_R n_12089 (.A1(n_11674_o_1),
    .A2(n_12073_o_0),
    .A3(n_12078_o_0),
    .B(n_12088_o_0),
    .Y(n_12089_o_0));
 NOR3xp33_ASAP7_75t_R n_1209 (.A(n_1006_o_0),
    .B(n_952_o_0),
    .C(n_878_o_0),
    .Y(n_1209_o_0));
 NAND2xp33_ASAP7_75t_R n_12090 (.A(n_11880_o_0),
    .B(n_11981_o_0),
    .Y(n_12090_o_0));
 OAI31xp33_ASAP7_75t_R n_12091 (.A1(n_11751_o_0),
    .A2(n_11764_o_0),
    .A3(n_11733_o_0),
    .B(n_11994_o_0),
    .Y(n_12091_o_0));
 AOI221xp5_ASAP7_75t_R n_12092 (.A1(n_11789_o_0),
    .A2(n_11840_o_0),
    .B1(n_11924_o_0),
    .B2(n_11923_o_0),
    .C(n_12091_o_0),
    .Y(n_12092_o_0));
 AOI31xp33_ASAP7_75t_R n_12093 (.A1(n_11763_o_0),
    .A2(n_12090_o_0),
    .A3(n_12043_o_0),
    .B(n_12092_o_0),
    .Y(n_12093_o_0));
 OAI21xp33_ASAP7_75t_R n_12094 (.A1(n_11766_o_0),
    .A2(n_11764_o_0),
    .B(n_11789_o_0),
    .Y(n_12094_o_0));
 AOI21xp33_ASAP7_75t_R n_12095 (.A1(n_11743_o_0),
    .A2(n_12094_o_0),
    .B(n_11896_o_0),
    .Y(n_12095_o_0));
 OAI31xp33_ASAP7_75t_R n_12096 (.A1(n_11796_o_0),
    .A2(n_11872_o_0),
    .A3(n_11918_o_0),
    .B(n_11798_o_0),
    .Y(n_12096_o_0));
 AOI21xp33_ASAP7_75t_R n_12097 (.A1(n_11845_o_0),
    .A2(n_12095_o_0),
    .B(n_12096_o_0),
    .Y(n_12097_o_0));
 AOI21xp33_ASAP7_75t_R n_12098 (.A1(n_11855_o_0),
    .A2(n_12097_o_0),
    .B(n_11675_o_0),
    .Y(n_12098_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_12099 (.A1(n_11764_o_0),
    .A2(n_11766_o_0),
    .B(n_11869_o_0),
    .C(n_11789_o_0),
    .D(n_11959_o_0),
    .Y(n_12099_o_0));
 AOI21xp33_ASAP7_75t_R n_1210 (.A1(n_1051_o_0),
    .A2(n_939_o_0),
    .B(n_904_o_0),
    .Y(n_1210_o_0));
 INVx1_ASAP7_75t_R n_12100 (.A(n_11881_o_0),
    .Y(n_12100_o_0));
 NAND3xp33_ASAP7_75t_R n_12101 (.A(n_11749_o_0),
    .B(n_11766_o_0),
    .C(n_11743_o_0),
    .Y(n_12101_o_0));
 OAI31xp33_ASAP7_75t_R n_12102 (.A1(n_11789_o_0),
    .A2(n_11787_o_0),
    .A3(n_12100_o_0),
    .B(n_12101_o_0),
    .Y(n_12102_o_0));
 OAI21xp33_ASAP7_75t_R n_12103 (.A1(n_11751_o_0),
    .A2(n_11843_o_0),
    .B(n_11761_o_0),
    .Y(n_12103_o_0));
 OAI21xp33_ASAP7_75t_R n_12104 (.A1(n_12074_o_0),
    .A2(n_12103_o_0),
    .B(n_11798_o_0),
    .Y(n_12104_o_0));
 OA211x2_ASAP7_75t_R n_12105 (.A1(n_11767_o_0),
    .A2(n_11766_o_0),
    .B(n_11751_o_0),
    .C(n_11811_o_0),
    .Y(n_12105_o_0));
 OAI21xp33_ASAP7_75t_R n_12106 (.A1(n_12105_o_0),
    .A2(n_12085_o_0),
    .B(n_11994_o_0),
    .Y(n_12106_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12107 (.A1(n_12102_o_0),
    .A2(n_11845_o_0),
    .B(n_12104_o_0),
    .C(n_12106_o_0),
    .Y(n_12107_o_0));
 AOI211xp5_ASAP7_75t_R n_12108 (.A1(n_12099_o_0),
    .A2(n_11754_o_0),
    .B(n_12107_o_0),
    .C(n_11674_o_1),
    .Y(n_12108_o_0));
 AOI211xp5_ASAP7_75t_R n_12109 (.A1(n_12093_o_0),
    .A2(n_12098_o_0),
    .B(n_12108_o_0),
    .C(n_11681_o_1),
    .Y(n_12109_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1211 (.A1(n_877_o_0),
    .A2(n_865_o_0),
    .B(n_1210_o_0),
    .C(n_891_o_0),
    .Y(n_1211_o_0));
 AOI21xp33_ASAP7_75t_R n_12110 (.A1(n_11857_o_0),
    .A2(n_12089_o_0),
    .B(n_12109_o_0),
    .Y(n_12110_o_0));
 AOI21xp33_ASAP7_75t_R n_12111 (.A1(n_11752_o_0),
    .A2(n_11751_o_0),
    .B(n_11745_o_0),
    .Y(n_12111_o_0));
 AOI221xp5_ASAP7_75t_R n_12112 (.A1(net76),
    .A2(n_11915_o_0),
    .B1(n_11766_o_0),
    .B2(n_11774_o_0),
    .C(n_11789_o_0),
    .Y(n_12112_o_0));
 AOI31xp33_ASAP7_75t_R n_12113 (.A1(n_11743_o_0),
    .A2(n_12023_o_0),
    .A3(n_11881_o_0),
    .B(n_12112_o_0),
    .Y(n_12113_o_0));
 OAI31xp33_ASAP7_75t_R n_12114 (.A1(n_11778_o_0),
    .A2(n_11852_o_0),
    .A3(n_11861_o_0),
    .B(n_11688_o_0),
    .Y(n_12114_o_0));
 AOI21xp33_ASAP7_75t_R n_12115 (.A1(n_12036_o_0),
    .A2(n_11767_o_0),
    .B(n_12114_o_0),
    .Y(n_12115_o_0));
 AOI21xp33_ASAP7_75t_R n_12116 (.A1(n_11798_o_0),
    .A2(n_12113_o_0),
    .B(n_12115_o_0),
    .Y(n_12116_o_0));
 NAND3xp33_ASAP7_75t_R n_12117 (.A(n_11817_o_0),
    .B(n_11805_o_0),
    .C(n_11789_o_0),
    .Y(n_12117_o_0));
 NAND2xp33_ASAP7_75t_R n_12118 (.A(n_11854_o_0),
    .B(n_11853_o_0),
    .Y(n_12118_o_0));
 AOI21xp33_ASAP7_75t_R n_12119 (.A1(n_12117_o_0),
    .A2(n_12118_o_0),
    .B(n_11959_o_0),
    .Y(n_12119_o_0));
 OAI21xp33_ASAP7_75t_R n_1212 (.A1(n_1208_o_0),
    .A2(n_1209_o_0),
    .B(n_1211_o_0),
    .Y(n_1212_o_0));
 AOI21xp33_ASAP7_75t_R n_12120 (.A1(n_11845_o_0),
    .A2(n_12116_o_0),
    .B(n_12119_o_0),
    .Y(n_12120_o_0));
 OAI21xp33_ASAP7_75t_R n_12121 (.A1(n_11965_o_0),
    .A2(n_12111_o_0),
    .B(n_12120_o_0),
    .Y(n_12121_o_0));
 OAI21xp33_ASAP7_75t_R n_12122 (.A1(n_11789_o_0),
    .A2(n_11803_o_0),
    .B(n_11688_o_0),
    .Y(n_12122_o_0));
 OAI21xp33_ASAP7_75t_R n_12123 (.A1(n_11789_o_0),
    .A2(n_12044_o_0),
    .B(n_11798_o_0),
    .Y(n_12123_o_0));
 AO21x1_ASAP7_75t_R n_12124 (.A1(n_11859_o_0),
    .A2(n_11941_o_0),
    .B(n_12123_o_0),
    .Y(n_12124_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12125 (.A1(n_11743_o_0),
    .A2(n_11941_o_0),
    .B(n_12122_o_0),
    .C(n_12124_o_0),
    .Y(n_12125_o_0));
 NOR2xp33_ASAP7_75t_R n_12126 (.A(n_1877_o_0),
    .B(n_11687_o_0),
    .Y(n_12126_o_0));
 AO21x1_ASAP7_75t_R n_12127 (.A1(n_11751_o_0),
    .A2(n_11880_o_0),
    .B(n_11836_o_0),
    .Y(n_12127_o_0));
 NAND2xp33_ASAP7_75t_R n_12128 (.A(n_11766_o_0),
    .B(n_11774_o_0),
    .Y(n_12128_o_0));
 OAI21xp33_ASAP7_75t_R n_12129 (.A1(n_11741_o_0),
    .A2(n_11777_o_0),
    .B(n_11733_o_0),
    .Y(n_12129_o_0));
 OAI31xp33_ASAP7_75t_R n_1213 (.A1(n_878_o_0),
    .A2(n_934_o_0),
    .A3(n_1088_o_0),
    .B(n_959_o_0),
    .Y(n_1213_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_12130 (.A1(n_11773_o_0),
    .A2(n_11824_o_0),
    .B(n_11884_o_0),
    .C(n_12129_o_0),
    .D(n_11861_o_0),
    .Y(n_12130_o_0));
 AOI31xp33_ASAP7_75t_R n_12131 (.A1(n_11751_o_0),
    .A2(n_12128_o_0),
    .A3(n_11809_o_0),
    .B(n_12130_o_0),
    .Y(n_12131_o_0));
 OAI21xp33_ASAP7_75t_R n_12132 (.A1(n_11798_o_0),
    .A2(n_12131_o_0),
    .B(n_11796_o_0),
    .Y(n_12132_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_12133 (.A1(n_1877_o_0),
    .A2(n_11687_o_0),
    .B(n_12126_o_0),
    .C(n_12127_o_0),
    .D(n_12132_o_0),
    .Y(n_12133_o_0));
 AOI211xp5_ASAP7_75t_R n_12134 (.A1(n_11782_o_0),
    .A2(n_12125_o_0),
    .B(n_12133_o_0),
    .C(n_11674_o_1),
    .Y(n_12134_o_0));
 AOI21xp33_ASAP7_75t_R n_12135 (.A1(n_11948_o_0),
    .A2(n_12121_o_0),
    .B(n_12134_o_0),
    .Y(n_12135_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12136 (.A1(net76),
    .A2(n_11752_o_0),
    .B(n_11766_o_0),
    .C(n_11924_o_0),
    .Y(n_12136_o_0));
 NAND2xp33_ASAP7_75t_R n_12137 (.A(n_11719_o_0),
    .B(n_12032_o_0),
    .Y(n_12137_o_0));
 OAI31xp33_ASAP7_75t_R n_12138 (.A1(n_11778_o_0),
    .A2(n_11787_o_0),
    .A3(n_11812_o_0),
    .B(n_12137_o_0),
    .Y(n_12138_o_0));
 AOI21xp33_ASAP7_75t_R n_12139 (.A1(n_11845_o_0),
    .A2(n_12138_o_0),
    .B(n_11675_o_0),
    .Y(n_12139_o_0));
 AOI21xp33_ASAP7_75t_R n_1214 (.A1(n_909_o_0),
    .A2(n_908_o_0),
    .B(n_903_o_0),
    .Y(n_1214_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12140 (.A1(n_11803_o_0),
    .A2(n_11733_o_0),
    .B(n_11852_o_0),
    .C(n_11778_o_0),
    .Y(n_12140_o_0));
 AOI31xp33_ASAP7_75t_R n_12141 (.A1(n_11743_o_0),
    .A2(n_11854_o_0),
    .A3(n_11892_o_0),
    .B(n_11761_o_0),
    .Y(n_12141_o_0));
 OAI21xp33_ASAP7_75t_R n_12142 (.A1(n_11789_o_0),
    .A2(n_11707_o_0),
    .B(n_12084_o_0),
    .Y(n_12142_o_0));
 AO21x1_ASAP7_75t_R n_12143 (.A1(n_12142_o_0),
    .A2(n_11761_o_0),
    .B(n_11948_o_0),
    .Y(n_12143_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12144 (.A1(n_12140_o_0),
    .A2(n_12141_o_0),
    .B(n_12143_o_0),
    .C(n_11689_o_0),
    .Y(n_12144_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_12145 (.A1(n_11841_o_0),
    .A2(n_12136_o_0),
    .B(n_11845_o_0),
    .C(n_12139_o_0),
    .D(n_12144_o_0),
    .Y(n_12145_o_0));
 OAI21xp33_ASAP7_75t_R n_12146 (.A1(n_11766_o_0),
    .A2(n_11913_o_0),
    .B(n_11918_o_0),
    .Y(n_12146_o_0));
 OAI32xp33_ASAP7_75t_R n_12147 (.A1(n_11845_o_0),
    .A2(n_12049_o_0),
    .A3(n_11779_o_0),
    .B1(n_12146_o_0),
    .B2(n_11761_o_0),
    .Y(n_12147_o_0));
 OAI32xp33_ASAP7_75t_R n_12148 (.A1(n_11743_o_0),
    .A2(n_11766_o_0),
    .A3(n_11774_o_0),
    .B1(n_12094_o_0),
    .B2(n_11956_o_0),
    .Y(n_12148_o_0));
 OAI21xp33_ASAP7_75t_R n_12149 (.A1(n_11778_o_0),
    .A2(n_11988_o_0),
    .B(n_11782_o_0),
    .Y(n_12149_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1215 (.A1(n_847_o_0),
    .A2(n_877_o_0),
    .B(n_1214_o_0),
    .C(net42),
    .Y(n_1215_o_0));
 AOI21xp33_ASAP7_75t_R n_12150 (.A1(n_11870_o_0),
    .A2(n_11916_o_0),
    .B(n_12149_o_0),
    .Y(n_12150_o_0));
 AOI211xp5_ASAP7_75t_R n_12151 (.A1(n_11796_o_0),
    .A2(n_12148_o_0),
    .B(n_12150_o_0),
    .C(n_11674_o_1),
    .Y(n_12151_o_0));
 AOI211xp5_ASAP7_75t_R n_12152 (.A1(n_11674_o_1),
    .A2(n_12147_o_0),
    .B(n_12151_o_0),
    .C(n_11798_o_0),
    .Y(n_12152_o_0));
 OAI22xp33_ASAP7_75t_R n_12153 (.A1(n_12145_o_0),
    .A2(n_12152_o_0),
    .B1(n_11829_o_0),
    .B2(n_11830_o_0),
    .Y(n_12153_o_0));
 OAI21xp33_ASAP7_75t_R n_12154 (.A1(n_11681_o_1),
    .A2(n_12135_o_0),
    .B(n_12153_o_0),
    .Y(n_12154_o_0));
 NAND2xp33_ASAP7_75t_R n_12155 (.A(n_11743_o_0),
    .B(n_11881_o_0),
    .Y(n_12155_o_0));
 INVx1_ASAP7_75t_R n_12156 (.A(n_12155_o_0),
    .Y(n_12156_o_0));
 AO21x1_ASAP7_75t_R n_12157 (.A1(n_11707_o_0),
    .A2(n_11766_o_0),
    .B(n_11906_o_0),
    .Y(n_12157_o_0));
 AOI22xp33_ASAP7_75t_R n_12158 (.A1(n_12156_o_0),
    .A2(n_12023_o_0),
    .B1(n_11751_o_0),
    .B2(n_12157_o_0),
    .Y(n_12158_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12159 (.A1(n_11766_o_0),
    .A2(n_11843_o_0),
    .B(n_11916_o_0),
    .C(n_11761_o_0),
    .Y(n_12159_o_0));
 OAI21xp33_ASAP7_75t_R n_1216 (.A1(n_904_o_0),
    .A2(n_1213_o_0),
    .B(n_1215_o_0),
    .Y(n_1216_o_0));
 AOI21xp33_ASAP7_75t_R n_12160 (.A1(n_11931_o_0),
    .A2(n_12159_o_0),
    .B(n_11799_o_0),
    .Y(n_12160_o_0));
 OAI21xp33_ASAP7_75t_R n_12161 (.A1(n_11848_o_0),
    .A2(n_11804_o_0),
    .B(n_11810_o_0),
    .Y(n_12161_o_0));
 OAI32xp33_ASAP7_75t_R n_12162 (.A1(n_11689_o_0),
    .A2(n_12161_o_0),
    .A3(n_11761_o_0),
    .B1(n_11959_o_0),
    .B2(n_11954_o_0),
    .Y(n_12162_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12163 (.A1(n_11796_o_0),
    .A2(n_12158_o_0),
    .B(n_12160_o_0),
    .C(n_12162_o_0),
    .Y(n_12163_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12164 (.A1(n_11999_o_0),
    .A2(n_11935_o_0),
    .B(n_11753_o_0),
    .C(n_11761_o_0),
    .Y(n_12164_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12165 (.A1(n_11751_o_0),
    .A2(n_11752_o_0),
    .B(net76),
    .C(n_11782_o_0),
    .Y(n_12165_o_0));
 AOI21xp33_ASAP7_75t_R n_12166 (.A1(n_11752_o_0),
    .A2(n_11733_o_0),
    .B(n_12165_o_0),
    .Y(n_12166_o_0));
 AO21x1_ASAP7_75t_R n_12167 (.A1(n_11859_o_0),
    .A2(n_11811_o_0),
    .B(n_11761_o_0),
    .Y(n_12167_o_0));
 AOI21xp33_ASAP7_75t_R n_12168 (.A1(n_11743_o_0),
    .A2(n_11895_o_0),
    .B(n_11845_o_0),
    .Y(n_12168_o_0));
 OAI21xp33_ASAP7_75t_R n_12169 (.A1(n_11915_o_0),
    .A2(n_11985_o_0),
    .B(n_11778_o_0),
    .Y(n_12169_o_0));
 NAND3xp33_ASAP7_75t_R n_1217 (.A(n_1212_o_0),
    .B(n_1216_o_0),
    .C(n_931_o_0),
    .Y(n_1217_o_0));
 AOI21xp33_ASAP7_75t_R n_12170 (.A1(n_12168_o_0),
    .A2(n_12169_o_0),
    .B(n_11798_o_0),
    .Y(n_12170_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12171 (.A1(n_11751_o_0),
    .A2(n_11793_o_0),
    .B(n_12167_o_0),
    .C(n_12170_o_0),
    .Y(n_12171_o_0));
 OAI31xp33_ASAP7_75t_R n_12172 (.A1(n_11688_o_0),
    .A2(n_12164_o_0),
    .A3(n_12166_o_0),
    .B(n_12171_o_0),
    .Y(n_12172_o_0));
 AOI22xp33_ASAP7_75t_R n_12173 (.A1(n_12163_o_0),
    .A2(n_11675_o_0),
    .B1(n_11948_o_0),
    .B2(n_12172_o_0),
    .Y(n_12173_o_0));
 OAI211xp5_ASAP7_75t_R n_12174 (.A1(n_11811_o_0),
    .A2(n_11707_o_0),
    .B(n_11751_o_0),
    .C(n_11753_o_0),
    .Y(n_12174_o_0));
 OAI31xp33_ASAP7_75t_R n_12175 (.A1(n_11778_o_0),
    .A2(n_11872_o_0),
    .A3(n_12044_o_0),
    .B(n_12174_o_0),
    .Y(n_12175_o_0));
 NAND3xp33_ASAP7_75t_R n_12176 (.A(n_11793_o_0),
    .B(n_11751_o_0),
    .C(n_11749_o_0),
    .Y(n_12176_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12177 (.A1(n_11803_o_0),
    .A2(n_12129_o_0),
    .B(n_12176_o_0),
    .C(n_11782_o_0),
    .Y(n_12177_o_0));
 AOI21xp33_ASAP7_75t_R n_12178 (.A1(n_11761_o_0),
    .A2(n_12175_o_0),
    .B(n_12177_o_0),
    .Y(n_12178_o_0));
 AOI311xp33_ASAP7_75t_R n_12179 (.A1(n_11766_o_0),
    .A2(n_11824_o_0),
    .A3(n_11773_o_0),
    .B(n_11778_o_0),
    .C(n_11869_o_0),
    .Y(n_12179_o_0));
 NAND2xp33_ASAP7_75t_R n_1218 (.A(n_836_o_0),
    .B(n_904_o_0),
    .Y(n_1218_o_0));
 AOI31xp33_ASAP7_75t_R n_12180 (.A1(n_11751_o_0),
    .A2(n_11927_o_0),
    .A3(n_11881_o_0),
    .B(n_12179_o_0),
    .Y(n_12180_o_0));
 OAI21xp33_ASAP7_75t_R n_12181 (.A1(n_11796_o_0),
    .A2(n_12180_o_0),
    .B(n_11798_o_0),
    .Y(n_12181_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12182 (.A1(n_11971_o_0),
    .A2(n_12056_o_0),
    .B(n_12181_o_0),
    .C(n_11675_o_0),
    .Y(n_12182_o_0));
 AOI21xp33_ASAP7_75t_R n_12183 (.A1(n_11688_o_0),
    .A2(n_12178_o_0),
    .B(n_12182_o_0),
    .Y(n_12183_o_0));
 NOR2xp33_ASAP7_75t_R n_12184 (.A(n_11733_o_0),
    .B(n_11767_o_0),
    .Y(n_12184_o_0));
 OAI21xp33_ASAP7_75t_R n_12185 (.A1(n_11752_o_0),
    .A2(n_11763_o_0),
    .B(n_11688_o_0),
    .Y(n_12185_o_0));
 AOI21xp33_ASAP7_75t_R n_12186 (.A1(n_11825_o_0),
    .A2(n_11981_o_0),
    .B(n_12185_o_0),
    .Y(n_12186_o_0));
 OAI21xp33_ASAP7_75t_R n_12187 (.A1(n_11930_o_0),
    .A2(n_11763_o_0),
    .B(n_11798_o_0),
    .Y(n_12187_o_0));
 AOI31xp33_ASAP7_75t_R n_12188 (.A1(n_11743_o_0),
    .A2(n_11766_o_0),
    .A3(n_11930_o_0),
    .B(n_12187_o_0),
    .Y(n_12188_o_0));
 OAI21xp33_ASAP7_75t_R n_12189 (.A1(n_12186_o_0),
    .A2(n_12188_o_0),
    .B(n_11796_o_0),
    .Y(n_12189_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1219 (.A1(n_935_o_0),
    .A2(n_1218_o_0),
    .B(n_1051_o_0),
    .C(n_829_o_0),
    .Y(n_1219_o_0));
 AOI21xp33_ASAP7_75t_R n_12190 (.A1(n_12184_o_0),
    .A2(n_11751_o_0),
    .B(n_12189_o_0),
    .Y(n_12190_o_0));
 OAI22xp33_ASAP7_75t_R n_12191 (.A1(n_11913_o_0),
    .A2(n_11984_o_0),
    .B1(n_11751_o_0),
    .B2(net76),
    .Y(n_12191_o_0));
 INVx1_ASAP7_75t_R n_12192 (.A(n_11935_o_0),
    .Y(n_12192_o_0));
 OAI211xp5_ASAP7_75t_R n_12193 (.A1(n_11764_o_0),
    .A2(n_11733_o_0),
    .B(n_11751_o_0),
    .C(n_11892_o_0),
    .Y(n_12193_o_0));
 OAI211xp5_ASAP7_75t_R n_12194 (.A1(n_12192_o_0),
    .A2(n_12070_o_0),
    .B(n_12193_o_0),
    .C(n_11782_o_0),
    .Y(n_12194_o_0));
 OAI32xp33_ASAP7_75t_R n_12195 (.A1(n_11845_o_0),
    .A2(n_11799_o_0),
    .A3(n_12191_o_0),
    .B1(n_12194_o_0),
    .B2(n_11689_o_0),
    .Y(n_12195_o_0));
 AOI211xp5_ASAP7_75t_R n_12196 (.A1(n_11674_o_0),
    .A2(n_11835_o_0),
    .B(n_12190_o_0),
    .C(n_12195_o_0),
    .Y(n_12196_o_0));
 OAI22xp33_ASAP7_75t_R n_12197 (.A1(n_12183_o_0),
    .A2(n_12196_o_0),
    .B1(n_11829_o_0),
    .B2(n_11830_o_0),
    .Y(n_12197_o_0));
 OAI21xp33_ASAP7_75t_R n_12198 (.A1(n_11681_o_1),
    .A2(n_12173_o_0),
    .B(n_12197_o_0),
    .Y(n_12198_o_0));
 AOI21xp33_ASAP7_75t_R n_12199 (.A1(n_11766_o_0),
    .A2(n_11930_o_0),
    .B(n_11840_o_0),
    .Y(n_12199_o_0));
 OAI21xp33_ASAP7_75t_R n_1220 (.A1(n_1061_o_0),
    .A2(n_917_o_0),
    .B(n_1219_o_0),
    .Y(n_1220_o_0));
 OAI21xp33_ASAP7_75t_R n_12200 (.A1(n_11787_o_0),
    .A2(n_11917_o_0),
    .B(n_11966_o_0),
    .Y(n_12200_o_0));
 OAI22xp33_ASAP7_75t_R n_12201 (.A1(n_11930_o_0),
    .A2(n_12129_o_0),
    .B1(n_11923_o_0),
    .B2(n_11789_o_0),
    .Y(n_12201_o_0));
 AOI21xp33_ASAP7_75t_R n_12202 (.A1(n_11766_o_0),
    .A2(n_11930_o_0),
    .B(n_12201_o_0),
    .Y(n_12202_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_12203 (.A1(n_11865_o_0),
    .A2(n_12199_o_0),
    .B(n_12200_o_0),
    .C(n_12202_o_0),
    .D(n_11959_o_0),
    .Y(n_12203_o_0));
 AOI211xp5_ASAP7_75t_R n_12204 (.A1(n_11865_o_0),
    .A2(n_12199_o_0),
    .B(n_12200_o_0),
    .C(n_12043_o_0),
    .Y(n_12204_o_0));
 AOI21xp33_ASAP7_75t_R n_12205 (.A1(n_11789_o_0),
    .A2(n_11863_o_0),
    .B(n_11798_o_0),
    .Y(n_12205_o_0));
 OAI21xp33_ASAP7_75t_R n_12206 (.A1(n_11787_o_0),
    .A2(n_11973_o_0),
    .B(n_11798_o_0),
    .Y(n_12206_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12207 (.A1(n_11892_o_0),
    .A2(n_12003_o_0),
    .B(n_12206_o_0),
    .C(n_11845_o_0),
    .Y(n_12207_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12208 (.A1(n_11913_o_0),
    .A2(n_11984_o_0),
    .B(n_12205_o_0),
    .C(n_12207_o_0),
    .Y(n_12208_o_0));
 NOR4xp25_ASAP7_75t_R n_12209 (.A(n_12203_o_0),
    .B(n_12204_o_0),
    .C(n_12208_o_0),
    .D(n_11675_o_0),
    .Y(n_12209_o_0));
 AOI31xp33_ASAP7_75t_R n_1221 (.A1(n_878_o_0),
    .A2(n_904_o_0),
    .A3(n_910_o_0),
    .B(n_1220_o_0),
    .Y(n_1221_o_0));
 INVx1_ASAP7_75t_R n_12210 (.A(n_12129_o_0),
    .Y(n_12210_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12211 (.A1(n_12210_o_0),
    .A2(n_11764_o_0),
    .B(n_11751_o_0),
    .C(n_11843_o_0),
    .Y(n_12211_o_0));
 OAI211xp5_ASAP7_75t_R n_12212 (.A1(n_11743_o_0),
    .A2(n_11940_o_0),
    .B(n_11837_o_0),
    .C(n_11799_o_0),
    .Y(n_12212_o_0));
 AOI31xp33_ASAP7_75t_R n_12213 (.A1(n_11774_o_0),
    .A2(n_11789_o_0),
    .A3(n_11733_o_0),
    .B(n_12212_o_0),
    .Y(n_12213_o_0));
 AOI211xp5_ASAP7_75t_R n_12214 (.A1(n_11798_o_0),
    .A2(n_12211_o_0),
    .B(n_12213_o_0),
    .C(n_11796_o_0),
    .Y(n_12214_o_0));
 NAND3xp33_ASAP7_75t_R n_12215 (.A(n_11793_o_0),
    .B(n_11749_o_0),
    .C(n_11743_o_0),
    .Y(n_12215_o_0));
 OAI22xp33_ASAP7_75t_R n_12216 (.A1(n_11895_o_0),
    .A2(n_11903_o_0),
    .B1(n_12155_o_0),
    .B2(n_11915_o_0),
    .Y(n_12216_o_0));
 OAI21xp33_ASAP7_75t_R n_12217 (.A1(n_11689_o_0),
    .A2(n_12216_o_0),
    .B(n_11845_o_0),
    .Y(n_12217_o_0));
 AOI21xp33_ASAP7_75t_R n_12218 (.A1(n_12215_o_0),
    .A2(n_11945_o_0),
    .B(n_12217_o_0),
    .Y(n_12218_o_0));
 NOR3xp33_ASAP7_75t_R n_12219 (.A(n_12214_o_0),
    .B(n_12218_o_0),
    .C(n_11948_o_0),
    .Y(n_12219_o_0));
 OAI211xp5_ASAP7_75t_R n_1222 (.A1(n_889_o_0),
    .A2(net32),
    .B(n_939_o_0),
    .C(n_877_o_0),
    .Y(n_1222_o_0));
 AOI31xp33_ASAP7_75t_R n_12220 (.A1(n_11743_o_0),
    .A2(n_11766_o_0),
    .A3(n_11774_o_0),
    .B(n_11845_o_0),
    .Y(n_12220_o_0));
 NAND3xp33_ASAP7_75t_R n_12221 (.A(n_11892_o_0),
    .B(n_11751_o_0),
    .C(n_11766_o_0),
    .Y(n_12221_o_0));
 OAI21xp33_ASAP7_75t_R n_12222 (.A1(n_11765_o_0),
    .A2(n_11794_o_0),
    .B(n_11796_o_0),
    .Y(n_12222_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12223 (.A1(n_11751_o_0),
    .A2(n_12076_o_0),
    .B(n_12222_o_0),
    .C(n_11799_o_0),
    .Y(n_12223_o_0));
 AOI21xp33_ASAP7_75t_R n_12224 (.A1(n_11719_o_0),
    .A2(n_11789_o_0),
    .B(n_12080_o_0),
    .Y(n_12224_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12225 (.A1(n_12155_o_0),
    .A2(n_11765_o_0),
    .B(n_12000_o_0),
    .C(n_11688_o_0),
    .Y(n_12225_o_0));
 OAI21xp33_ASAP7_75t_R n_12226 (.A1(n_11761_o_0),
    .A2(n_12224_o_0),
    .B(n_12225_o_0),
    .Y(n_12226_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12227 (.A1(n_12220_o_0),
    .A2(n_12221_o_0),
    .B(n_12223_o_0),
    .C(n_12226_o_0),
    .Y(n_12227_o_0));
 INVx1_ASAP7_75t_R n_12228 (.A(n_11844_o_0),
    .Y(n_12228_o_0));
 AOI22xp33_ASAP7_75t_R n_12229 (.A1(n_12156_o_0),
    .A2(n_11719_o_0),
    .B1(n_12228_o_0),
    .B2(n_12199_o_0),
    .Y(n_12229_o_0));
 OAI31xp33_ASAP7_75t_R n_1223 (.A1(n_1050_o_0),
    .A2(n_1146_o_0),
    .A3(n_877_o_0),
    .B(n_1222_o_0),
    .Y(n_1223_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_12230 (.A1(n_11848_o_0),
    .A2(n_11804_o_0),
    .B(n_12192_o_0),
    .C(n_11845_o_0),
    .Y(n_12230_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12231 (.A1(n_11796_o_0),
    .A2(n_12229_o_0),
    .B(n_12230_o_0),
    .C(n_11798_o_0),
    .Y(n_12231_o_0));
 OAI21xp33_ASAP7_75t_R n_12232 (.A1(n_12070_o_0),
    .A2(n_12192_o_0),
    .B(n_12009_o_0),
    .Y(n_12232_o_0));
 AOI31xp33_ASAP7_75t_R n_12233 (.A1(n_11796_o_0),
    .A2(n_11904_o_0),
    .A3(n_12059_o_0),
    .B(n_11689_o_0),
    .Y(n_12233_o_0));
 OAI21xp33_ASAP7_75t_R n_12234 (.A1(n_11796_o_0),
    .A2(n_12232_o_0),
    .B(n_12233_o_0),
    .Y(n_12234_o_0));
 AOI31xp33_ASAP7_75t_R n_12235 (.A1(n_11948_o_0),
    .A2(n_12231_o_0),
    .A3(n_12234_o_0),
    .B(n_11857_o_0),
    .Y(n_12235_o_0));
 OAI21xp33_ASAP7_75t_R n_12236 (.A1(n_11948_o_0),
    .A2(n_12227_o_0),
    .B(n_12235_o_0),
    .Y(n_12236_o_0));
 OAI31xp33_ASAP7_75t_R n_12237 (.A1(n_11831_o_0),
    .A2(n_12209_o_0),
    .A3(n_12219_o_0),
    .B(n_12236_o_0),
    .Y(n_12237_o_0));
 INVx1_ASAP7_75t_R n_12238 (.A(_00645_),
    .Y(n_12238_o_0));
 INVx1_ASAP7_75t_R n_12239 (.A(_00647_),
    .Y(n_12239_o_0));
 AOI21xp33_ASAP7_75t_R n_1224 (.A1(n_877_o_0),
    .A2(n_984_o_0),
    .B(n_1121_o_0),
    .Y(n_1224_o_0));
 INVx1_ASAP7_75t_R n_12240 (.A(_00729_),
    .Y(n_12240_o_0));
 NOR5xp2_ASAP7_75t_R n_12241 (.A(n_12238_o_0),
    .B(n_12239_o_0),
    .C(n_12240_o_0),
    .D(ld),
    .E(_00648_),
    .Y(n_12241_o_0));
 XOR2xp5_ASAP7_75t_R n_12242 (.A(_00860_),
    .B(_01115_),
    .Y(n_12242_o_0));
 XOR2xp5_ASAP7_75t_R n_12243 (.A(_00861_),
    .B(_01116_),
    .Y(n_12243_o_0));
 XOR2xp5_ASAP7_75t_R n_12244 (.A(_00862_),
    .B(_01117_),
    .Y(n_12244_o_0));
 XOR2xp5_ASAP7_75t_R n_12245 (.A(_00863_),
    .B(_01118_),
    .Y(n_12245_o_0));
 XOR2xp5_ASAP7_75t_R n_12246 (.A(_00864_),
    .B(_01119_),
    .Y(n_12246_o_0));
 XOR2xp5_ASAP7_75t_R n_12247 (.A(_00865_),
    .B(_01120_),
    .Y(n_12247_o_0));
 XOR2xp5_ASAP7_75t_R n_12248 (.A(_00866_),
    .B(_01121_),
    .Y(n_12248_o_0));
 XOR2xp5_ASAP7_75t_R n_12249 (.A(_00642_),
    .B(_00867_),
    .Y(n_12249_o_0));
 AOI21xp33_ASAP7_75t_R n_1225 (.A1(net42),
    .A2(n_1224_o_0),
    .B(n_903_o_0),
    .Y(n_1225_o_0));
 XOR2xp5_ASAP7_75t_R n_12250 (.A(_00868_),
    .B(_01076_),
    .Y(n_12250_o_0));
 XOR2xp5_ASAP7_75t_R n_12251 (.A(_00869_),
    .B(_01077_),
    .Y(n_12251_o_0));
 XOR2xp5_ASAP7_75t_R n_12252 (.A(_00870_),
    .B(_01078_),
    .Y(n_12252_o_0));
 XOR2xp5_ASAP7_75t_R n_12253 (.A(_00871_),
    .B(_01079_),
    .Y(n_12253_o_0));
 XOR2xp5_ASAP7_75t_R n_12254 (.A(_00872_),
    .B(_01080_),
    .Y(n_12254_o_0));
 XOR2xp5_ASAP7_75t_R n_12255 (.A(_00873_),
    .B(_01081_),
    .Y(n_12255_o_0));
 XOR2xp5_ASAP7_75t_R n_12256 (.A(_00874_),
    .B(_01082_),
    .Y(n_12256_o_0));
 XOR2xp5_ASAP7_75t_R n_12257 (.A(_00643_),
    .B(_00875_),
    .Y(n_12257_o_0));
 XOR2xp5_ASAP7_75t_R n_12258 (.A(_00876_),
    .B(_01036_),
    .Y(n_12258_o_0));
 XOR2xp5_ASAP7_75t_R n_12259 (.A(_00877_),
    .B(_01037_),
    .Y(n_12259_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1226 (.A1(net15),
    .A2(n_1223_o_0),
    .B(n_903_o_0),
    .C(n_1225_o_0),
    .Y(n_1226_o_0));
 XOR2xp5_ASAP7_75t_R n_12260 (.A(_00878_),
    .B(_01038_),
    .Y(n_12260_o_0));
 XOR2xp5_ASAP7_75t_R n_12261 (.A(_00879_),
    .B(_01039_),
    .Y(n_12261_o_0));
 XOR2xp5_ASAP7_75t_R n_12262 (.A(_00880_),
    .B(_01040_),
    .Y(n_12262_o_0));
 XOR2xp5_ASAP7_75t_R n_12263 (.A(_00881_),
    .B(_01041_),
    .Y(n_12263_o_0));
 XOR2xp5_ASAP7_75t_R n_12264 (.A(_00882_),
    .B(_01042_),
    .Y(n_12264_o_0));
 XOR2xp5_ASAP7_75t_R n_12265 (.A(_00883_),
    .B(_01043_),
    .Y(n_12265_o_0));
 XOR2xp5_ASAP7_75t_R n_12266 (.A(_00884_),
    .B(_00996_),
    .Y(n_12266_o_0));
 XOR2xp5_ASAP7_75t_R n_12267 (.A(_00885_),
    .B(_00997_),
    .Y(n_12267_o_0));
 XOR2xp5_ASAP7_75t_R n_12268 (.A(_00886_),
    .B(_00998_),
    .Y(n_12268_o_0));
 XOR2xp5_ASAP7_75t_R n_12269 (.A(_00887_),
    .B(_00999_),
    .Y(n_12269_o_0));
 OAI21xp33_ASAP7_75t_R n_1227 (.A1(n_1221_o_0),
    .A2(n_1226_o_0),
    .B(n_930_o_0),
    .Y(n_1227_o_0));
 XOR2xp5_ASAP7_75t_R n_12270 (.A(_00888_),
    .B(_01000_),
    .Y(n_12270_o_0));
 XOR2xp5_ASAP7_75t_R n_12271 (.A(_00889_),
    .B(_01001_),
    .Y(n_12271_o_0));
 XOR2xp5_ASAP7_75t_R n_12272 (.A(_00890_),
    .B(_01002_),
    .Y(n_12272_o_0));
 XOR2xp5_ASAP7_75t_R n_12273 (.A(_00891_),
    .B(_01003_),
    .Y(n_12273_o_0));
 XOR2xp5_ASAP7_75t_R n_12274 (.A(_00964_),
    .B(_01068_),
    .Y(n_12274_o_0));
 XOR2xp5_ASAP7_75t_R n_12275 (.A(_00965_),
    .B(_01069_),
    .Y(n_12275_o_0));
 XOR2xp5_ASAP7_75t_R n_12276 (.A(_00966_),
    .B(_01070_),
    .Y(n_12276_o_0));
 XOR2xp5_ASAP7_75t_R n_12277 (.A(_00967_),
    .B(_01071_),
    .Y(n_12277_o_0));
 XOR2xp5_ASAP7_75t_R n_12278 (.A(_00968_),
    .B(_01072_),
    .Y(n_12278_o_0));
 XOR2xp5_ASAP7_75t_R n_12279 (.A(_00969_),
    .B(_01073_),
    .Y(n_12279_o_0));
 OAI21xp33_ASAP7_75t_R n_1228 (.A1(n_972_o_0),
    .A2(n_1217_o_0),
    .B(n_1227_o_0),
    .Y(n_1228_o_0));
 XOR2xp5_ASAP7_75t_R n_12280 (.A(_00970_),
    .B(_01074_),
    .Y(n_12280_o_0));
 XOR2xp5_ASAP7_75t_R n_12281 (.A(_00971_),
    .B(_01075_),
    .Y(n_12281_o_0));
 XOR2xp5_ASAP7_75t_R n_12282 (.A(_00972_),
    .B(_01028_),
    .Y(n_12282_o_0));
 XOR2xp5_ASAP7_75t_R n_12283 (.A(_00973_),
    .B(_01029_),
    .Y(n_12283_o_0));
 XOR2xp5_ASAP7_75t_R n_12284 (.A(_00974_),
    .B(_01030_),
    .Y(n_12284_o_0));
 XOR2xp5_ASAP7_75t_R n_12285 (.A(_00975_),
    .B(_01031_),
    .Y(n_12285_o_0));
 XOR2xp5_ASAP7_75t_R n_12286 (.A(_00976_),
    .B(_01032_),
    .Y(n_12286_o_0));
 XOR2xp5_ASAP7_75t_R n_12287 (.A(_00977_),
    .B(_01033_),
    .Y(n_12287_o_0));
 XOR2xp5_ASAP7_75t_R n_12288 (.A(_00978_),
    .B(_01034_),
    .Y(n_12288_o_0));
 XOR2xp5_ASAP7_75t_R n_12289 (.A(_00979_),
    .B(_01035_),
    .Y(n_12289_o_0));
 NOR2xp33_ASAP7_75t_R n_1229 (.A(n_859_o_0),
    .B(net32),
    .Y(n_1229_o_0));
 XOR2xp5_ASAP7_75t_R n_12290 (.A(_00980_),
    .B(_01020_),
    .Y(n_12290_o_0));
 XOR2xp5_ASAP7_75t_R n_12291 (.A(_00981_),
    .B(_01021_),
    .Y(n_12291_o_0));
 XOR2xp5_ASAP7_75t_R n_12292 (.A(_00982_),
    .B(_01022_),
    .Y(n_12292_o_0));
 XOR2xp5_ASAP7_75t_R n_12293 (.A(_00983_),
    .B(_01023_),
    .Y(n_12293_o_0));
 XOR2xp5_ASAP7_75t_R n_12294 (.A(_00984_),
    .B(_01024_),
    .Y(n_12294_o_0));
 XOR2xp5_ASAP7_75t_R n_12295 (.A(_00985_),
    .B(_01025_),
    .Y(n_12295_o_0));
 XOR2xp5_ASAP7_75t_R n_12296 (.A(_00986_),
    .B(_01026_),
    .Y(n_12296_o_0));
 XOR2xp5_ASAP7_75t_R n_12297 (.A(_00987_),
    .B(_01027_),
    .Y(n_12297_o_0));
 XOR2xp5_ASAP7_75t_R n_12298 (.A(_00924_),
    .B(_01099_),
    .Y(n_12298_o_0));
 XOR2xp5_ASAP7_75t_R n_12299 (.A(_00925_),
    .B(_01100_),
    .Y(n_12299_o_0));
 OAI31xp33_ASAP7_75t_R n_1230 (.A1(n_878_o_0),
    .A2(n_915_o_0),
    .A3(n_1229_o_0),
    .B(n_1045_o_0),
    .Y(n_1230_o_0));
 XOR2xp5_ASAP7_75t_R n_12300 (.A(_00926_),
    .B(_01101_),
    .Y(n_12300_o_0));
 XOR2xp5_ASAP7_75t_R n_12301 (.A(_00927_),
    .B(_01102_),
    .Y(n_12301_o_0));
 XOR2xp5_ASAP7_75t_R n_12302 (.A(_00928_),
    .B(_01103_),
    .Y(n_12302_o_0));
 XOR2xp5_ASAP7_75t_R n_12303 (.A(_00929_),
    .B(_01104_),
    .Y(n_12303_o_0));
 XOR2xp5_ASAP7_75t_R n_12304 (.A(_00930_),
    .B(_01105_),
    .Y(n_12304_o_0));
 XOR2xp5_ASAP7_75t_R n_12305 (.A(_00931_),
    .B(_01106_),
    .Y(n_12305_o_0));
 XOR2xp5_ASAP7_75t_R n_12306 (.A(_00932_),
    .B(_01060_),
    .Y(n_12306_o_0));
 XOR2xp5_ASAP7_75t_R n_12307 (.A(_00933_),
    .B(_01061_),
    .Y(n_12307_o_0));
 XOR2xp5_ASAP7_75t_R n_12308 (.A(_00934_),
    .B(_01062_),
    .Y(n_12308_o_0));
 XOR2xp5_ASAP7_75t_R n_12309 (.A(_00935_),
    .B(_01063_),
    .Y(n_12309_o_0));
 OAI21xp33_ASAP7_75t_R n_1231 (.A1(n_881_o_0),
    .A2(n_957_o_0),
    .B(n_877_o_0),
    .Y(n_1231_o_0));
 XOR2xp5_ASAP7_75t_R n_12310 (.A(_00936_),
    .B(_01064_),
    .Y(n_12310_o_0));
 XOR2xp5_ASAP7_75t_R n_12311 (.A(_00937_),
    .B(_01065_),
    .Y(n_12311_o_0));
 XOR2xp5_ASAP7_75t_R n_12312 (.A(_00938_),
    .B(_01066_),
    .Y(n_12312_o_0));
 XOR2xp5_ASAP7_75t_R n_12313 (.A(_00939_),
    .B(_01067_),
    .Y(n_12313_o_0));
 XOR2xp5_ASAP7_75t_R n_12314 (.A(_00940_),
    .B(_01052_),
    .Y(n_12314_o_0));
 XOR2xp5_ASAP7_75t_R n_12315 (.A(_00941_),
    .B(_01053_),
    .Y(n_12315_o_0));
 XOR2xp5_ASAP7_75t_R n_12316 (.A(_00942_),
    .B(_01054_),
    .Y(n_12316_o_0));
 XOR2xp5_ASAP7_75t_R n_12317 (.A(_00943_),
    .B(_01055_),
    .Y(n_12317_o_0));
 XOR2xp5_ASAP7_75t_R n_12318 (.A(_00944_),
    .B(_01056_),
    .Y(n_12318_o_0));
 XOR2xp5_ASAP7_75t_R n_12319 (.A(_00945_),
    .B(_01057_),
    .Y(n_12319_o_0));
 OAI21xp33_ASAP7_75t_R n_1232 (.A1(n_915_o_0),
    .A2(n_883_o_0),
    .B(n_1231_o_0),
    .Y(n_1232_o_0));
 XOR2xp5_ASAP7_75t_R n_12320 (.A(_00946_),
    .B(_01058_),
    .Y(n_12320_o_0));
 XOR2xp5_ASAP7_75t_R n_12321 (.A(_00947_),
    .B(_01059_),
    .Y(n_12321_o_0));
 XOR2xp5_ASAP7_75t_R n_12322 (.A(_00948_),
    .B(_01012_),
    .Y(n_12322_o_0));
 XOR2xp5_ASAP7_75t_R n_12323 (.A(_00949_),
    .B(_01013_),
    .Y(n_12323_o_0));
 XOR2xp5_ASAP7_75t_R n_12324 (.A(_00950_),
    .B(_01014_),
    .Y(n_12324_o_0));
 XOR2xp5_ASAP7_75t_R n_12325 (.A(_00951_),
    .B(_01015_),
    .Y(n_12325_o_0));
 XOR2xp5_ASAP7_75t_R n_12326 (.A(_00952_),
    .B(_01016_),
    .Y(n_12326_o_0));
 XOR2xp5_ASAP7_75t_R n_12327 (.A(_00953_),
    .B(_01017_),
    .Y(n_12327_o_0));
 XOR2xp5_ASAP7_75t_R n_12328 (.A(_00954_),
    .B(_01018_),
    .Y(n_12328_o_0));
 XOR2xp5_ASAP7_75t_R n_12329 (.A(_00955_),
    .B(_01019_),
    .Y(n_12329_o_0));
 OAI21xp33_ASAP7_75t_R n_1233 (.A1(net42),
    .A2(n_1232_o_0),
    .B(n_903_o_0),
    .Y(n_1233_o_0));
 XOR2xp5_ASAP7_75t_R n_12330 (.A(_00892_),
    .B(_01091_),
    .Y(n_12330_o_0));
 XOR2xp5_ASAP7_75t_R n_12331 (.A(_00893_),
    .B(_01092_),
    .Y(n_12331_o_0));
 XOR2xp5_ASAP7_75t_R n_12332 (.A(_00894_),
    .B(_01093_),
    .Y(n_12332_o_0));
 XOR2xp5_ASAP7_75t_R n_12333 (.A(_00895_),
    .B(_01094_),
    .Y(n_12333_o_0));
 XOR2xp5_ASAP7_75t_R n_12334 (.A(_00896_),
    .B(_01095_),
    .Y(n_12334_o_0));
 XOR2xp5_ASAP7_75t_R n_12335 (.A(_00897_),
    .B(_01096_),
    .Y(n_12335_o_0));
 XOR2xp5_ASAP7_75t_R n_12336 (.A(_00898_),
    .B(_01097_),
    .Y(n_12336_o_0));
 XOR2xp5_ASAP7_75t_R n_12337 (.A(_00899_),
    .B(_01098_),
    .Y(n_12337_o_0));
 XOR2xp5_ASAP7_75t_R n_12338 (.A(_00900_),
    .B(_01083_),
    .Y(n_12338_o_0));
 XOR2xp5_ASAP7_75t_R n_12339 (.A(_00901_),
    .B(_01084_),
    .Y(n_12339_o_0));
 NAND2xp33_ASAP7_75t_R n_1234 (.A(n_933_o_0),
    .B(n_877_o_0),
    .Y(n_1234_o_0));
 XOR2xp5_ASAP7_75t_R n_12340 (.A(_00902_),
    .B(_01085_),
    .Y(n_12340_o_0));
 XOR2xp5_ASAP7_75t_R n_12341 (.A(_00903_),
    .B(_01086_),
    .Y(n_12341_o_0));
 XOR2xp5_ASAP7_75t_R n_12342 (.A(_00904_),
    .B(_01087_),
    .Y(n_12342_o_0));
 XOR2xp5_ASAP7_75t_R n_12343 (.A(_00905_),
    .B(_01088_),
    .Y(n_12343_o_0));
 XOR2xp5_ASAP7_75t_R n_12344 (.A(_00906_),
    .B(_01089_),
    .Y(n_12344_o_0));
 XOR2xp5_ASAP7_75t_R n_12345 (.A(_00907_),
    .B(_01090_),
    .Y(n_12345_o_0));
 XOR2xp5_ASAP7_75t_R n_12346 (.A(_00956_),
    .B(_01107_),
    .Y(n_12346_o_0));
 XOR2xp5_ASAP7_75t_R n_12347 (.A(_00957_),
    .B(_01108_),
    .Y(n_12347_o_0));
 XOR2xp5_ASAP7_75t_R n_12348 (.A(_00958_),
    .B(_01109_),
    .Y(n_12348_o_0));
 XOR2xp5_ASAP7_75t_R n_12349 (.A(_00959_),
    .B(_01110_),
    .Y(n_12349_o_0));
 AOI21xp33_ASAP7_75t_R n_1235 (.A1(n_1234_o_0),
    .A2(n_864_o_0),
    .B(n_1190_o_0),
    .Y(n_1235_o_0));
 XOR2xp5_ASAP7_75t_R n_12350 (.A(_00960_),
    .B(_01111_),
    .Y(n_12350_o_0));
 XOR2xp5_ASAP7_75t_R n_12351 (.A(_00961_),
    .B(_01112_),
    .Y(n_12351_o_0));
 XOR2xp5_ASAP7_75t_R n_12352 (.A(_00962_),
    .B(_01113_),
    .Y(n_12352_o_0));
 XOR2xp5_ASAP7_75t_R n_12353 (.A(_00963_),
    .B(_01114_),
    .Y(n_12353_o_0));
 XOR2xp5_ASAP7_75t_R n_12354 (.A(_00908_),
    .B(_01044_),
    .Y(n_12354_o_0));
 XOR2xp5_ASAP7_75t_R n_12355 (.A(_00909_),
    .B(_01045_),
    .Y(n_12355_o_0));
 XOR2xp5_ASAP7_75t_R n_12356 (.A(_00910_),
    .B(_01046_),
    .Y(n_12356_o_0));
 XOR2xp5_ASAP7_75t_R n_12357 (.A(_00911_),
    .B(_01047_),
    .Y(n_12357_o_0));
 XOR2xp5_ASAP7_75t_R n_12358 (.A(_00912_),
    .B(_01048_),
    .Y(n_12358_o_0));
 XOR2xp5_ASAP7_75t_R n_12359 (.A(_00913_),
    .B(_01049_),
    .Y(n_12359_o_0));
 OAI211xp5_ASAP7_75t_R n_1236 (.A1(n_913_o_0),
    .A2(n_836_o_0),
    .B(n_865_o_0),
    .C(n_878_o_0),
    .Y(n_1236_o_0));
 XOR2xp5_ASAP7_75t_R n_12360 (.A(_00914_),
    .B(_01050_),
    .Y(n_12360_o_0));
 XOR2xp5_ASAP7_75t_R n_12361 (.A(_00915_),
    .B(_01051_),
    .Y(n_12361_o_0));
 XOR2xp5_ASAP7_75t_R n_12362 (.A(_00916_),
    .B(_01004_),
    .Y(n_12362_o_0));
 XOR2xp5_ASAP7_75t_R n_12363 (.A(_00917_),
    .B(_01005_),
    .Y(n_12363_o_0));
 XOR2xp5_ASAP7_75t_R n_12364 (.A(_00918_),
    .B(_01006_),
    .Y(n_12364_o_0));
 XOR2xp5_ASAP7_75t_R n_12365 (.A(_00919_),
    .B(_01007_),
    .Y(n_12365_o_0));
 XOR2xp5_ASAP7_75t_R n_12366 (.A(_00920_),
    .B(_01008_),
    .Y(n_12366_o_0));
 XOR2xp5_ASAP7_75t_R n_12367 (.A(_00921_),
    .B(_01009_),
    .Y(n_12367_o_0));
 XOR2xp5_ASAP7_75t_R n_12368 (.A(_00922_),
    .B(_01010_),
    .Y(n_12368_o_0));
 XOR2xp5_ASAP7_75t_R n_12369 (.A(_00923_),
    .B(_01011_),
    .Y(n_12369_o_0));
 OAI211xp5_ASAP7_75t_R n_1237 (.A1(n_847_o_0),
    .A2(n_859_o_0),
    .B(n_944_o_0),
    .C(n_877_o_0),
    .Y(n_1237_o_0));
 NAND2xp33_ASAP7_75t_R n_12370 (.A(key[96]),
    .B(ld),
    .Y(n_12370_o_0));
 OAI21xp33_ASAP7_75t_R n_12371 (.A1(ld),
    .A2(n_1900_o_0),
    .B(n_12370_o_0),
    .Y(n_12371_o_0));
 INVx1_ASAP7_75t_R n_12372 (.A(key[106]),
    .Y(n_12372_o_0));
 AOI21xp33_ASAP7_75t_R n_12373 (.A1(n_12372_o_0),
    .A2(ld),
    .B(n_1366_o_0),
    .Y(n_12373_o_0));
 INVx1_ASAP7_75t_R n_12374 (.A(n_1392_o_0),
    .Y(n_12374_o_0));
 NAND2xp33_ASAP7_75t_R n_12375 (.A(key[107]),
    .B(ld),
    .Y(n_12375_o_0));
 OAI21xp33_ASAP7_75t_R n_12376 (.A1(ld),
    .A2(n_12374_o_0),
    .B(n_12375_o_0),
    .Y(n_12376_o_0));
 INVx1_ASAP7_75t_R n_12377 (.A(n_1356_o_0),
    .Y(n_12377_o_0));
 NAND2xp33_ASAP7_75t_R n_12378 (.A(key[108]),
    .B(ld),
    .Y(n_12378_o_0));
 OAI21xp33_ASAP7_75t_R n_12379 (.A1(ld),
    .A2(n_12377_o_0),
    .B(n_12378_o_0),
    .Y(n_12379_o_0));
 AOI31xp33_ASAP7_75t_R n_1238 (.A1(net42),
    .A2(n_1236_o_0),
    .A3(n_1237_o_0),
    .B(n_903_o_0),
    .Y(n_1238_o_0));
 INVx1_ASAP7_75t_R n_12380 (.A(n_1419_o_0),
    .Y(n_12380_o_0));
 NAND2xp33_ASAP7_75t_R n_12381 (.A(key[109]),
    .B(ld),
    .Y(n_12381_o_0));
 OAI21xp33_ASAP7_75t_R n_12382 (.A1(ld),
    .A2(n_12380_o_0),
    .B(n_12381_o_0),
    .Y(n_12382_o_0));
 NAND2xp33_ASAP7_75t_R n_12383 (.A(key[110]),
    .B(ld),
    .Y(n_12383_o_0));
 OAI21xp33_ASAP7_75t_R n_12384 (.A1(ld),
    .A2(n_1348_o_0),
    .B(n_12383_o_0),
    .Y(n_12384_o_0));
 NAND2xp33_ASAP7_75t_R n_12385 (.A(key[111]),
    .B(ld),
    .Y(n_12385_o_0));
 OAI21xp33_ASAP7_75t_R n_12386 (.A1(ld),
    .A2(n_1339_o_0),
    .B(n_12385_o_0),
    .Y(n_12386_o_0));
 INVx1_ASAP7_75t_R n_12387 (.A(n_838_o_0),
    .Y(n_12387_o_0));
 NAND2xp33_ASAP7_75t_R n_12388 (.A(key[112]),
    .B(ld),
    .Y(n_12388_o_0));
 OAI21xp33_ASAP7_75t_R n_12389 (.A1(ld),
    .A2(n_12387_o_0),
    .B(n_12388_o_0),
    .Y(n_12389_o_0));
 OAI21xp33_ASAP7_75t_R n_1239 (.A1(net42),
    .A2(n_1235_o_0),
    .B(n_1238_o_0),
    .Y(n_1239_o_0));
 INVx1_ASAP7_75t_R n_12390 (.A(n_850_o_0),
    .Y(n_12390_o_0));
 NAND2xp33_ASAP7_75t_R n_12391 (.A(key[113]),
    .B(ld),
    .Y(n_12391_o_0));
 OAI21xp33_ASAP7_75t_R n_12392 (.A1(ld),
    .A2(n_12390_o_0),
    .B(n_12391_o_0),
    .Y(n_12392_o_0));
 NAND2xp33_ASAP7_75t_R n_12393 (.A(key[114]),
    .B(ld),
    .Y(n_12393_o_0));
 OAI21xp33_ASAP7_75t_R n_12394 (.A1(ld),
    .A2(n_832_o_0),
    .B(n_12393_o_0),
    .Y(n_12394_o_0));
 INVx1_ASAP7_75t_R n_12395 (.A(n_867_o_0),
    .Y(n_12395_o_0));
 NAND2xp33_ASAP7_75t_R n_12396 (.A(key[115]),
    .B(ld),
    .Y(n_12396_o_0));
 OAI21xp33_ASAP7_75t_R n_12397 (.A1(ld),
    .A2(n_12395_o_0),
    .B(n_12396_o_0),
    .Y(n_12397_o_0));
 NAND2xp33_ASAP7_75t_R n_12398 (.A(key[97]),
    .B(ld),
    .Y(n_12398_o_0));
 OAI21xp33_ASAP7_75t_R n_12399 (.A1(ld),
    .A2(n_1905_o_0),
    .B(n_12398_o_0),
    .Y(n_12399_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1240 (.A1(net16),
    .A2(n_1230_o_0),
    .B(n_1233_o_0),
    .C(n_1239_o_0),
    .Y(n_1240_o_0));
 INVx1_ASAP7_75t_R n_12400 (.A(n_822_o_0),
    .Y(n_12400_o_0));
 NAND2xp33_ASAP7_75t_R n_12401 (.A(key[116]),
    .B(ld),
    .Y(n_12401_o_0));
 OAI21xp33_ASAP7_75t_R n_12402 (.A1(ld),
    .A2(n_12400_o_0),
    .B(n_12401_o_0),
    .Y(n_12402_o_0));
 INVx1_ASAP7_75t_R n_12403 (.A(n_895_o_0),
    .Y(n_12403_o_0));
 NAND2xp33_ASAP7_75t_R n_12404 (.A(key[117]),
    .B(ld),
    .Y(n_12404_o_0));
 OAI21xp33_ASAP7_75t_R n_12405 (.A1(ld),
    .A2(n_12403_o_0),
    .B(n_12404_o_0),
    .Y(n_12405_o_0));
 NAND2xp33_ASAP7_75t_R n_12406 (.A(key[118]),
    .B(ld),
    .Y(n_12406_o_0));
 OAI21xp33_ASAP7_75t_R n_12407 (.A1(ld),
    .A2(n_924_o_0),
    .B(n_12406_o_0),
    .Y(n_12407_o_0));
 NAND2xp33_ASAP7_75t_R n_12408 (.A(key[119]),
    .B(ld),
    .Y(n_12408_o_0));
 OAI21xp33_ASAP7_75t_R n_12409 (.A1(ld),
    .A2(n_965_o_0),
    .B(n_12408_o_0),
    .Y(n_12409_o_0));
 AOI21xp33_ASAP7_75t_R n_1241 (.A1(n_877_o_0),
    .A2(n_882_o_0),
    .B(net16),
    .Y(n_1241_o_0));
 NAND2xp33_ASAP7_75t_R n_12410 (.A(key[120]),
    .B(ld),
    .Y(n_12410_o_0));
 OAI21xp33_ASAP7_75t_R n_12411 (.A1(ld),
    .A2(n_2493_o_0),
    .B(n_12410_o_0),
    .Y(n_12411_o_0));
 NAND2xp33_ASAP7_75t_R n_12412 (.A(key[121]),
    .B(ld),
    .Y(n_12412_o_0));
 OAI21xp33_ASAP7_75t_R n_12413 (.A1(ld),
    .A2(n_2454_o_0),
    .B(n_12412_o_0),
    .Y(n_12413_o_0));
 NAND2xp33_ASAP7_75t_R n_12414 (.A(key[122]),
    .B(ld),
    .Y(n_12414_o_0));
 OAI31xp33_ASAP7_75t_R n_12415 (.A1(ld),
    .A2(n_2479_o_0),
    .A3(n_2477_o_0),
    .B(n_12414_o_0),
    .Y(n_12415_o_0));
 NAND2xp33_ASAP7_75t_R n_12416 (.A(key[123]),
    .B(ld),
    .Y(n_12416_o_0));
 OAI21xp33_ASAP7_75t_R n_12417 (.A1(ld),
    .A2(n_2408_o_0),
    .B(n_12416_o_0),
    .Y(n_12417_o_0));
 NAND2xp33_ASAP7_75t_R n_12418 (.A(key[124]),
    .B(ld),
    .Y(n_12418_o_0));
 OAI21xp33_ASAP7_75t_R n_12419 (.A1(ld),
    .A2(n_2517_o_0),
    .B(n_12418_o_0),
    .Y(n_12419_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1242 (.A1(n_881_o_0),
    .A2(n_935_o_0),
    .B(n_878_o_0),
    .C(n_829_o_0),
    .Y(n_1242_o_0));
 INVx1_ASAP7_75t_R n_12420 (.A(n_2388_o_0),
    .Y(n_12420_o_0));
 NAND2xp33_ASAP7_75t_R n_12421 (.A(key[125]),
    .B(ld),
    .Y(n_12421_o_0));
 OAI21xp33_ASAP7_75t_R n_12422 (.A1(ld),
    .A2(n_12420_o_0),
    .B(n_12421_o_0),
    .Y(n_12422_o_0));
 INVx1_ASAP7_75t_R n_12423 (.A(key[98]),
    .Y(n_12423_o_0));
 AOI21xp33_ASAP7_75t_R n_12424 (.A1(n_12423_o_0),
    .A2(ld),
    .B(n_1892_o_0),
    .Y(n_12424_o_0));
 INVx1_ASAP7_75t_R n_12425 (.A(n_2376_o_0),
    .Y(n_12425_o_0));
 NAND2xp33_ASAP7_75t_R n_12426 (.A(key[126]),
    .B(ld),
    .Y(n_12426_o_0));
 OAI21xp33_ASAP7_75t_R n_12427 (.A1(ld),
    .A2(n_12425_o_0),
    .B(n_12426_o_0),
    .Y(n_12427_o_0));
 NAND2xp33_ASAP7_75t_R n_12428 (.A(key[127]),
    .B(ld),
    .Y(n_12428_o_0));
 OAI21xp33_ASAP7_75t_R n_12429 (.A1(ld),
    .A2(n_2365_o_0),
    .B(n_12428_o_0),
    .Y(n_12429_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1243 (.A1(n_935_o_0),
    .A2(net32),
    .B(n_1242_o_0),
    .C(n_903_o_0),
    .Y(n_1243_o_0));
 INVx1_ASAP7_75t_R n_12430 (.A(n_1919_o_0),
    .Y(n_12430_o_0));
 NAND2xp33_ASAP7_75t_R n_12431 (.A(key[99]),
    .B(ld),
    .Y(n_12431_o_0));
 OAI21xp33_ASAP7_75t_R n_12432 (.A1(ld),
    .A2(n_12430_o_0),
    .B(n_12431_o_0),
    .Y(n_12432_o_0));
 INVx1_ASAP7_75t_R n_12433 (.A(n_1881_o_0),
    .Y(n_12433_o_0));
 NAND2xp33_ASAP7_75t_R n_12434 (.A(key[100]),
    .B(ld),
    .Y(n_12434_o_0));
 OAI21xp33_ASAP7_75t_R n_12435 (.A1(ld),
    .A2(n_12433_o_0),
    .B(n_12434_o_0),
    .Y(n_12435_o_0));
 INVx1_ASAP7_75t_R n_12436 (.A(n_1874_o_0),
    .Y(n_12436_o_0));
 NAND2xp33_ASAP7_75t_R n_12437 (.A(key[101]),
    .B(ld),
    .Y(n_12437_o_0));
 OAI21xp33_ASAP7_75t_R n_12438 (.A1(ld),
    .A2(n_12436_o_0),
    .B(n_12437_o_0),
    .Y(n_12438_o_0));
 NAND2xp33_ASAP7_75t_R n_12439 (.A(key[102]),
    .B(ld),
    .Y(n_12439_o_0));
 AOI21xp33_ASAP7_75t_R n_1244 (.A1(n_1156_o_0),
    .A2(n_1241_o_0),
    .B(n_1243_o_0),
    .Y(n_1244_o_0));
 OAI21xp33_ASAP7_75t_R n_12440 (.A1(ld),
    .A2(n_1866_o_0),
    .B(n_12439_o_0),
    .Y(n_12440_o_0));
 NAND2xp33_ASAP7_75t_R n_12441 (.A(key[103]),
    .B(ld),
    .Y(n_12441_o_0));
 OAI21xp33_ASAP7_75t_R n_12442 (.A1(ld),
    .A2(n_1859_o_0),
    .B(n_12441_o_0),
    .Y(n_12442_o_0));
 NAND2xp33_ASAP7_75t_R n_12443 (.A(key[104]),
    .B(ld),
    .Y(n_12443_o_0));
 OAI21xp33_ASAP7_75t_R n_12444 (.A1(ld),
    .A2(n_1382_o_0),
    .B(n_12443_o_0),
    .Y(n_12444_o_0));
 NAND2xp33_ASAP7_75t_R n_12445 (.A(key[105]),
    .B(ld),
    .Y(n_12445_o_0));
 OAI21xp33_ASAP7_75t_R n_12446 (.A1(ld),
    .A2(n_1373_o_0),
    .B(n_12445_o_0),
    .Y(n_12446_o_0));
 NAND2xp33_ASAP7_75t_R n_12447 (.A(key[64]),
    .B(ld),
    .Y(n_12447_o_0));
 OAI21xp33_ASAP7_75t_R n_12448 (.A1(ld),
    .A2(n_1902_o_0),
    .B(n_12447_o_0),
    .Y(n_12448_o_0));
 NAND2xp33_ASAP7_75t_R n_12449 (.A(n_8305_o_0),
    .B(n_1365_o_0),
    .Y(n_12449_o_0));
 OAI21xp33_ASAP7_75t_R n_1245 (.A1(n_1190_o_0),
    .A2(n_1121_o_0),
    .B(n_941_o_0),
    .Y(n_1245_o_0));
 OAI21xp33_ASAP7_75t_R n_12450 (.A1(n_1365_o_0),
    .A2(n_8305_o_0),
    .B(n_12449_o_0),
    .Y(n_12450_o_0));
 NAND2xp33_ASAP7_75t_R n_12451 (.A(key[74]),
    .B(ld),
    .Y(n_12451_o_0));
 OAI21xp33_ASAP7_75t_R n_12452 (.A1(ld),
    .A2(n_12450_o_0),
    .B(n_12451_o_0),
    .Y(n_12452_o_0));
 NAND2xp33_ASAP7_75t_R n_12453 (.A(key[75]),
    .B(ld),
    .Y(n_12453_o_0));
 OAI21xp33_ASAP7_75t_R n_12454 (.A1(ld),
    .A2(n_1395_o_0),
    .B(n_12453_o_0),
    .Y(n_12454_o_0));
 INVx1_ASAP7_75t_R n_12455 (.A(n_1357_o_0),
    .Y(n_12455_o_0));
 NAND2xp33_ASAP7_75t_R n_12456 (.A(key[76]),
    .B(ld),
    .Y(n_12456_o_0));
 OAI21xp33_ASAP7_75t_R n_12457 (.A1(ld),
    .A2(n_12455_o_0),
    .B(n_12456_o_0),
    .Y(n_12457_o_0));
 INVx1_ASAP7_75t_R n_12458 (.A(n_1420_o_0),
    .Y(n_12458_o_0));
 NAND2xp33_ASAP7_75t_R n_12459 (.A(key[77]),
    .B(ld),
    .Y(n_12459_o_0));
 INVx1_ASAP7_75t_R n_1246 (.A(n_995_o_0),
    .Y(n_1246_o_0));
 OAI21xp33_ASAP7_75t_R n_12460 (.A1(ld),
    .A2(n_12458_o_0),
    .B(n_12459_o_0),
    .Y(n_12460_o_0));
 NAND2xp33_ASAP7_75t_R n_12461 (.A(key[78]),
    .B(ld),
    .Y(n_12461_o_0));
 OAI21xp33_ASAP7_75t_R n_12462 (.A1(ld),
    .A2(n_1350_o_0),
    .B(n_12461_o_0),
    .Y(n_12462_o_0));
 INVx1_ASAP7_75t_R n_12463 (.A(n_1341_o_0),
    .Y(n_12463_o_0));
 NAND2xp33_ASAP7_75t_R n_12464 (.A(key[79]),
    .B(ld),
    .Y(n_12464_o_0));
 OAI21xp33_ASAP7_75t_R n_12465 (.A1(ld),
    .A2(n_12463_o_0),
    .B(n_12464_o_0),
    .Y(n_12465_o_0));
 NAND2xp33_ASAP7_75t_R n_12466 (.A(key[80]),
    .B(ld),
    .Y(n_12466_o_0));
 OAI21xp33_ASAP7_75t_R n_12467 (.A1(ld),
    .A2(n_841_o_0),
    .B(n_12466_o_0),
    .Y(n_12467_o_0));
 NAND2xp33_ASAP7_75t_R n_12468 (.A(key[81]),
    .B(ld),
    .Y(n_12468_o_0));
 OAI21xp33_ASAP7_75t_R n_12469 (.A1(ld),
    .A2(n_855_o_0),
    .B(n_12468_o_0),
    .Y(n_12469_o_0));
 OAI31xp33_ASAP7_75t_R n_1247 (.A1(n_877_o_0),
    .A2(n_1088_o_0),
    .A3(n_907_o_0),
    .B(n_829_o_0),
    .Y(n_1247_o_0));
 XNOR2xp5_ASAP7_75t_R n_12470 (.A(_00910_),
    .B(n_832_o_0),
    .Y(n_12470_o_0));
 NAND2xp33_ASAP7_75t_R n_12471 (.A(key[82]),
    .B(ld),
    .Y(n_12471_o_0));
 OAI21xp33_ASAP7_75t_R n_12472 (.A1(ld),
    .A2(n_12470_o_0),
    .B(n_12471_o_0),
    .Y(n_12472_o_0));
 NAND2xp33_ASAP7_75t_R n_12473 (.A(key[83]),
    .B(ld),
    .Y(n_12473_o_0));
 OAI21xp33_ASAP7_75t_R n_12474 (.A1(ld),
    .A2(n_870_o_0),
    .B(n_12473_o_0),
    .Y(n_12474_o_0));
 NAND2xp33_ASAP7_75t_R n_12475 (.A(key[65]),
    .B(ld),
    .Y(n_12475_o_0));
 OAI21xp33_ASAP7_75t_R n_12476 (.A1(ld),
    .A2(n_1907_o_0),
    .B(n_12475_o_0),
    .Y(n_12476_o_0));
 INVx1_ASAP7_75t_R n_12477 (.A(n_823_o_0),
    .Y(n_12477_o_0));
 NAND2xp33_ASAP7_75t_R n_12478 (.A(key[84]),
    .B(ld),
    .Y(n_12478_o_0));
 OAI21xp33_ASAP7_75t_R n_12479 (.A1(ld),
    .A2(n_12477_o_0),
    .B(n_12478_o_0),
    .Y(n_12479_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1248 (.A1(n_1246_o_0),
    .A2(n_1005_o_0),
    .B(n_1247_o_0),
    .C(n_904_o_0),
    .Y(n_1248_o_0));
 NAND2xp33_ASAP7_75t_R n_12480 (.A(key[85]),
    .B(ld),
    .Y(n_12480_o_0));
 OAI21xp33_ASAP7_75t_R n_12481 (.A1(ld),
    .A2(n_896_o_0),
    .B(n_12480_o_0),
    .Y(n_12481_o_0));
 NAND2xp33_ASAP7_75t_R n_12482 (.A(key[86]),
    .B(ld),
    .Y(n_12482_o_0));
 OAI21xp33_ASAP7_75t_R n_12483 (.A1(ld),
    .A2(n_925_o_0),
    .B(n_12482_o_0),
    .Y(n_12483_o_0));
 NAND2xp33_ASAP7_75t_R n_12484 (.A(key[87]),
    .B(ld),
    .Y(n_12484_o_0));
 OAI21xp33_ASAP7_75t_R n_12485 (.A1(ld),
    .A2(n_966_o_0),
    .B(n_12484_o_0),
    .Y(n_12485_o_0));
 NAND2xp33_ASAP7_75t_R n_12486 (.A(key[88]),
    .B(ld),
    .Y(n_12486_o_0));
 OAI31xp33_ASAP7_75t_R n_12487 (.A1(ld),
    .A2(n_2425_o_0),
    .A3(n_2422_o_0),
    .B(n_12486_o_0),
    .Y(n_12487_o_0));
 NAND2xp33_ASAP7_75t_R n_12488 (.A(key[89]),
    .B(ld),
    .Y(n_12488_o_0));
 OAI31xp33_ASAP7_75t_R n_12489 (.A1(ld),
    .A2(n_2443_o_0),
    .A3(n_2501_o_0),
    .B(n_12488_o_0),
    .Y(n_12489_o_0));
 AOI21xp33_ASAP7_75t_R n_1249 (.A1(n_960_o_0),
    .A2(n_1245_o_0),
    .B(n_1248_o_0),
    .Y(n_1249_o_0));
 NAND2xp33_ASAP7_75t_R n_12490 (.A(key[90]),
    .B(ld),
    .Y(n_12490_o_0));
 OAI31xp33_ASAP7_75t_R n_12491 (.A1(ld),
    .A2(n_2489_o_0),
    .A3(n_2472_o_0),
    .B(n_12490_o_0),
    .Y(n_12491_o_0));
 AND2x2_ASAP7_75t_R n_12492 (.A(key[91]),
    .B(ld),
    .Y(n_12492_o_0));
 AOI31xp33_ASAP7_75t_R n_12493 (.A1(n_827_o_0),
    .A2(n_2405_o_0),
    .A3(n_2401_o_0),
    .B(n_12492_o_0),
    .Y(n_12493_o_0));
 INVx1_ASAP7_75t_R n_12494 (.A(n_12493_o_0),
    .Y(n_12494_o_0));
 INVx1_ASAP7_75t_R n_12495 (.A(n_2519_o_0),
    .Y(n_12495_o_0));
 NAND2xp33_ASAP7_75t_R n_12496 (.A(key[92]),
    .B(ld),
    .Y(n_12496_o_0));
 OAI21xp33_ASAP7_75t_R n_12497 (.A1(ld),
    .A2(n_12495_o_0),
    .B(n_12496_o_0),
    .Y(n_12497_o_0));
 INVx1_ASAP7_75t_R n_12498 (.A(n_2389_o_0),
    .Y(n_12498_o_0));
 NAND2xp33_ASAP7_75t_R n_12499 (.A(key[93]),
    .B(ld),
    .Y(n_12499_o_0));
 OAI21xp33_ASAP7_75t_R n_1250 (.A1(n_1244_o_0),
    .A2(n_1249_o_0),
    .B(n_931_o_0),
    .Y(n_1250_o_0));
 OAI21xp33_ASAP7_75t_R n_12500 (.A1(ld),
    .A2(n_12498_o_0),
    .B(n_12499_o_0),
    .Y(n_12500_o_0));
 NAND2xp33_ASAP7_75t_R n_12501 (.A(_00894_),
    .B(n_1891_o_0),
    .Y(n_12501_o_0));
 OAI21xp33_ASAP7_75t_R n_12502 (.A1(_00894_),
    .A2(n_1891_o_0),
    .B(n_12501_o_0),
    .Y(n_12502_o_0));
 NAND2xp33_ASAP7_75t_R n_12503 (.A(key[66]),
    .B(ld),
    .Y(n_12503_o_0));
 OAI21xp33_ASAP7_75t_R n_12504 (.A1(ld),
    .A2(n_12502_o_0),
    .B(n_12503_o_0),
    .Y(n_12504_o_0));
 INVx1_ASAP7_75t_R n_12505 (.A(n_2377_o_0),
    .Y(n_12505_o_0));
 NAND2xp33_ASAP7_75t_R n_12506 (.A(key[94]),
    .B(ld),
    .Y(n_12506_o_0));
 OAI21xp33_ASAP7_75t_R n_12507 (.A1(ld),
    .A2(n_12505_o_0),
    .B(n_12506_o_0),
    .Y(n_12507_o_0));
 NAND2xp33_ASAP7_75t_R n_12508 (.A(key[95]),
    .B(ld),
    .Y(n_12508_o_0));
 OAI21xp33_ASAP7_75t_R n_12509 (.A1(ld),
    .A2(n_2366_o_0),
    .B(n_12508_o_0),
    .Y(n_12509_o_0));
 OAI21xp33_ASAP7_75t_R n_1251 (.A1(n_931_o_0),
    .A2(n_1240_o_0),
    .B(n_1250_o_0),
    .Y(n_1251_o_0));
 INVx1_ASAP7_75t_R n_12510 (.A(n_1920_o_0),
    .Y(n_12510_o_0));
 NAND2xp33_ASAP7_75t_R n_12511 (.A(key[67]),
    .B(ld),
    .Y(n_12511_o_0));
 OAI21xp33_ASAP7_75t_R n_12512 (.A1(ld),
    .A2(n_12510_o_0),
    .B(n_12511_o_0),
    .Y(n_12512_o_0));
 INVx1_ASAP7_75t_R n_12513 (.A(n_1882_o_0),
    .Y(n_12513_o_0));
 NAND2xp33_ASAP7_75t_R n_12514 (.A(key[68]),
    .B(ld),
    .Y(n_12514_o_0));
 OAI21xp33_ASAP7_75t_R n_12515 (.A1(ld),
    .A2(n_12513_o_0),
    .B(n_12514_o_0),
    .Y(n_12515_o_0));
 INVx1_ASAP7_75t_R n_12516 (.A(n_1875_o_0),
    .Y(n_12516_o_0));
 NAND2xp33_ASAP7_75t_R n_12517 (.A(key[69]),
    .B(ld),
    .Y(n_12517_o_0));
 OAI21xp33_ASAP7_75t_R n_12518 (.A1(ld),
    .A2(n_12516_o_0),
    .B(n_12517_o_0),
    .Y(n_12518_o_0));
 NAND2xp33_ASAP7_75t_R n_12519 (.A(key[70]),
    .B(ld),
    .Y(n_12519_o_0));
 NAND2xp33_ASAP7_75t_R n_1252 (.A(n_972_o_0),
    .B(n_1251_o_0),
    .Y(n_1252_o_0));
 OAI21xp33_ASAP7_75t_R n_12520 (.A1(ld),
    .A2(n_1867_o_0),
    .B(n_12519_o_0),
    .Y(n_12520_o_0));
 NAND2xp33_ASAP7_75t_R n_12521 (.A(key[71]),
    .B(ld),
    .Y(n_12521_o_0));
 OAI21xp33_ASAP7_75t_R n_12522 (.A1(ld),
    .A2(n_1860_o_0),
    .B(n_12521_o_0),
    .Y(n_12522_o_0));
 NAND2xp33_ASAP7_75t_R n_12523 (.A(key[72]),
    .B(ld),
    .Y(n_12523_o_0));
 OAI21xp33_ASAP7_75t_R n_12524 (.A1(ld),
    .A2(n_1384_o_0),
    .B(n_12523_o_0),
    .Y(n_12524_o_0));
 NAND2xp33_ASAP7_75t_R n_12525 (.A(key[73]),
    .B(ld),
    .Y(n_12525_o_0));
 OAI21xp33_ASAP7_75t_R n_12526 (.A1(ld),
    .A2(n_1375_o_0),
    .B(n_12525_o_0),
    .Y(n_12526_o_0));
 XNOR2xp5_ASAP7_75t_R n_12527 (.A(_00924_),
    .B(n_1902_o_0),
    .Y(n_12527_o_0));
 NAND2xp33_ASAP7_75t_R n_12528 (.A(key[32]),
    .B(ld),
    .Y(n_12528_o_0));
 OAI21xp33_ASAP7_75t_R n_12529 (.A1(ld),
    .A2(n_12527_o_0),
    .B(n_12528_o_0),
    .Y(n_12529_o_0));
 OAI21xp33_ASAP7_75t_R n_1253 (.A1(n_972_o_0),
    .A2(n_1228_o_0),
    .B(n_1252_o_0),
    .Y(n_1253_o_0));
 XNOR2xp5_ASAP7_75t_R n_12530 (.A(_00934_),
    .B(n_12450_o_0),
    .Y(n_12530_o_0));
 NAND2xp33_ASAP7_75t_R n_12531 (.A(key[42]),
    .B(ld),
    .Y(n_12531_o_0));
 OAI21xp33_ASAP7_75t_R n_12532 (.A1(ld),
    .A2(n_12530_o_0),
    .B(n_12531_o_0),
    .Y(n_12532_o_0));
 XNOR2xp5_ASAP7_75t_R n_12533 (.A(_00935_),
    .B(n_1395_o_0),
    .Y(n_12533_o_0));
 NAND2xp33_ASAP7_75t_R n_12534 (.A(key[43]),
    .B(ld),
    .Y(n_12534_o_0));
 OAI21xp33_ASAP7_75t_R n_12535 (.A1(ld),
    .A2(n_12533_o_0),
    .B(n_12534_o_0),
    .Y(n_12535_o_0));
 INVx1_ASAP7_75t_R n_12536 (.A(n_1358_o_0),
    .Y(n_12536_o_0));
 NAND2xp33_ASAP7_75t_R n_12537 (.A(key[44]),
    .B(ld),
    .Y(n_12537_o_0));
 OAI21xp33_ASAP7_75t_R n_12538 (.A1(ld),
    .A2(n_12536_o_0),
    .B(n_12537_o_0),
    .Y(n_12538_o_0));
 NAND2xp33_ASAP7_75t_R n_12539 (.A(key[45]),
    .B(ld),
    .Y(n_12539_o_0));
 NAND3xp33_ASAP7_75t_R n_1254 (.A(n_993_o_0),
    .B(n_909_o_0),
    .C(n_878_o_0),
    .Y(n_1254_o_0));
 OAI21xp33_ASAP7_75t_R n_12540 (.A1(ld),
    .A2(n_1493_o_0),
    .B(n_12539_o_0),
    .Y(n_12540_o_0));
 NAND2xp33_ASAP7_75t_R n_12541 (.A(key[46]),
    .B(ld),
    .Y(n_12541_o_0));
 OAI21xp33_ASAP7_75t_R n_12542 (.A1(ld),
    .A2(n_1352_o_0),
    .B(n_12541_o_0),
    .Y(n_12542_o_0));
 NAND2xp33_ASAP7_75t_R n_12543 (.A(key[47]),
    .B(ld),
    .Y(n_12543_o_0));
 OAI21xp33_ASAP7_75t_R n_12544 (.A1(ld),
    .A2(n_1344_o_0),
    .B(n_12543_o_0),
    .Y(n_12544_o_0));
 XNOR2xp5_ASAP7_75t_R n_12545 (.A(_00940_),
    .B(n_841_o_0),
    .Y(n_12545_o_0));
 NAND2xp33_ASAP7_75t_R n_12546 (.A(key[48]),
    .B(ld),
    .Y(n_12546_o_0));
 OAI21xp33_ASAP7_75t_R n_12547 (.A1(ld),
    .A2(n_12545_o_0),
    .B(n_12546_o_0),
    .Y(n_12547_o_0));
 XNOR2xp5_ASAP7_75t_R n_12548 (.A(_00941_),
    .B(n_855_o_0),
    .Y(n_12548_o_0));
 NAND2xp33_ASAP7_75t_R n_12549 (.A(key[49]),
    .B(ld),
    .Y(n_12549_o_0));
 OAI31xp33_ASAP7_75t_R n_1255 (.A1(n_878_o_0),
    .A2(n_952_o_0),
    .A3(n_1088_o_0),
    .B(n_1254_o_0),
    .Y(n_1255_o_0));
 OAI21xp33_ASAP7_75t_R n_12550 (.A1(ld),
    .A2(n_12548_o_0),
    .B(n_12549_o_0),
    .Y(n_12550_o_0));
 XNOR2xp5_ASAP7_75t_R n_12551 (.A(_00942_),
    .B(n_12470_o_0),
    .Y(n_12551_o_0));
 NAND2xp33_ASAP7_75t_R n_12552 (.A(key[50]),
    .B(ld),
    .Y(n_12552_o_0));
 OAI21xp33_ASAP7_75t_R n_12553 (.A1(ld),
    .A2(n_12551_o_0),
    .B(n_12552_o_0),
    .Y(n_12553_o_0));
 AOI211xp5_ASAP7_75t_R n_12554 (.A1(n_870_o_0),
    .A2(_00943_),
    .B(n_871_o_0),
    .C(ld),
    .Y(n_12554_o_0));
 AO21x1_ASAP7_75t_R n_12555 (.A1(key[51]),
    .A2(ld),
    .B(n_12554_o_0),
    .Y(n_12555_o_0));
 XNOR2xp5_ASAP7_75t_R n_12556 (.A(_00925_),
    .B(n_1907_o_0),
    .Y(n_12556_o_0));
 NAND2xp33_ASAP7_75t_R n_12557 (.A(key[33]),
    .B(ld),
    .Y(n_12557_o_0));
 OAI21xp33_ASAP7_75t_R n_12558 (.A1(ld),
    .A2(n_12556_o_0),
    .B(n_12557_o_0),
    .Y(n_12558_o_0));
 INVx1_ASAP7_75t_R n_12559 (.A(n_824_o_0),
    .Y(n_12559_o_0));
 AOI21xp33_ASAP7_75t_R n_1256 (.A1(n_1167_o_0),
    .A2(n_1254_o_0),
    .B(n_994_o_0),
    .Y(n_1256_o_0));
 NAND2xp33_ASAP7_75t_R n_12560 (.A(key[52]),
    .B(ld),
    .Y(n_12560_o_0));
 OAI21xp33_ASAP7_75t_R n_12561 (.A1(ld),
    .A2(n_12559_o_0),
    .B(n_12560_o_0),
    .Y(n_12561_o_0));
 AOI211xp5_ASAP7_75t_R n_12562 (.A1(n_896_o_0),
    .A2(_00945_),
    .B(n_897_o_0),
    .C(ld),
    .Y(n_12562_o_0));
 AO21x1_ASAP7_75t_R n_12563 (.A1(key[53]),
    .A2(ld),
    .B(n_12562_o_0),
    .Y(n_12563_o_0));
 INVx1_ASAP7_75t_R n_12564 (.A(n_927_o_0),
    .Y(n_12564_o_0));
 NAND2xp33_ASAP7_75t_R n_12565 (.A(key[54]),
    .B(ld),
    .Y(n_12565_o_0));
 OAI21xp33_ASAP7_75t_R n_12566 (.A1(ld),
    .A2(n_12564_o_0),
    .B(n_12565_o_0),
    .Y(n_12566_o_0));
 NAND2xp33_ASAP7_75t_R n_12567 (.A(key[55]),
    .B(ld),
    .Y(n_12567_o_0));
 OAI21xp33_ASAP7_75t_R n_12568 (.A1(ld),
    .A2(n_967_o_0),
    .B(n_12567_o_0),
    .Y(n_12568_o_0));
 NAND2xp33_ASAP7_75t_R n_12569 (.A(key[56]),
    .B(ld),
    .Y(n_12569_o_0));
 OAI21xp33_ASAP7_75t_R n_1257 (.A1(n_903_o_0),
    .A2(n_1256_o_0),
    .B(net16),
    .Y(n_1257_o_0));
 OAI31xp33_ASAP7_75t_R n_12570 (.A1(ld),
    .A2(n_2494_o_0),
    .A3(n_2434_o_0),
    .B(n_12569_o_0),
    .Y(n_12570_o_0));
 INVx1_ASAP7_75t_R n_12571 (.A(n_2536_o_0),
    .Y(n_12571_o_0));
 NAND2xp33_ASAP7_75t_R n_12572 (.A(key[57]),
    .B(ld),
    .Y(n_12572_o_0));
 OAI21xp33_ASAP7_75t_R n_12573 (.A1(ld),
    .A2(n_12571_o_0),
    .B(n_12572_o_0),
    .Y(n_12573_o_0));
 INVx1_ASAP7_75t_R n_12574 (.A(n_2476_o_0),
    .Y(n_12574_o_0));
 NAND2xp33_ASAP7_75t_R n_12575 (.A(key[58]),
    .B(ld),
    .Y(n_12575_o_0));
 OAI21xp33_ASAP7_75t_R n_12576 (.A1(ld),
    .A2(n_12574_o_0),
    .B(n_12575_o_0),
    .Y(n_12576_o_0));
 INVx1_ASAP7_75t_R n_12577 (.A(n_2409_o_0),
    .Y(n_12577_o_0));
 NAND2xp33_ASAP7_75t_R n_12578 (.A(key[59]),
    .B(ld),
    .Y(n_12578_o_0));
 OAI31xp33_ASAP7_75t_R n_12579 (.A1(ld),
    .A2(n_12577_o_0),
    .A3(n_2412_o_0),
    .B(n_12578_o_0),
    .Y(n_12579_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1258 (.A1(n_904_o_0),
    .A2(n_1255_o_0),
    .B(net16),
    .C(n_1257_o_0),
    .Y(n_1258_o_0));
 INVx1_ASAP7_75t_R n_12580 (.A(n_2522_o_0),
    .Y(n_12580_o_0));
 NAND2xp33_ASAP7_75t_R n_12581 (.A(key[60]),
    .B(ld),
    .Y(n_12581_o_0));
 OAI31xp33_ASAP7_75t_R n_12582 (.A1(ld),
    .A2(n_12580_o_0),
    .A3(n_2524_o_0),
    .B(n_12581_o_0),
    .Y(n_12582_o_0));
 INVx1_ASAP7_75t_R n_12583 (.A(n_2529_o_0),
    .Y(n_12583_o_0));
 NAND2xp33_ASAP7_75t_R n_12584 (.A(key[61]),
    .B(ld),
    .Y(n_12584_o_0));
 OAI21xp33_ASAP7_75t_R n_12585 (.A1(ld),
    .A2(n_12583_o_0),
    .B(n_12584_o_0),
    .Y(n_12585_o_0));
 XNOR2xp5_ASAP7_75t_R n_12586 (.A(_00926_),
    .B(n_12502_o_0),
    .Y(n_12586_o_0));
 NAND2xp33_ASAP7_75t_R n_12587 (.A(key[34]),
    .B(ld),
    .Y(n_12587_o_0));
 OAI21xp33_ASAP7_75t_R n_12588 (.A1(ld),
    .A2(n_12586_o_0),
    .B(n_12587_o_0),
    .Y(n_12588_o_0));
 NAND2xp33_ASAP7_75t_R n_12589 (.A(key[62]),
    .B(ld),
    .Y(n_12589_o_0));
 OAI21xp33_ASAP7_75t_R n_1259 (.A1(n_934_o_0),
    .A2(n_936_o_0),
    .B(net16),
    .Y(n_1259_o_0));
 OAI21xp33_ASAP7_75t_R n_12590 (.A1(ld),
    .A2(n_2380_o_0),
    .B(n_12589_o_0),
    .Y(n_12590_o_0));
 INVx1_ASAP7_75t_R n_12591 (.A(n_2368_o_0),
    .Y(n_12591_o_0));
 NAND2xp33_ASAP7_75t_R n_12592 (.A(key[63]),
    .B(ld),
    .Y(n_12592_o_0));
 OAI21xp33_ASAP7_75t_R n_12593 (.A1(ld),
    .A2(n_12591_o_0),
    .B(n_12592_o_0),
    .Y(n_12593_o_0));
 INVx1_ASAP7_75t_R n_12594 (.A(n_1921_o_0),
    .Y(n_12594_o_0));
 NAND2xp33_ASAP7_75t_R n_12595 (.A(key[35]),
    .B(ld),
    .Y(n_12595_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_12596 (.A1(n_12594_o_0),
    .A2(n_1924_o_0),
    .B(ld),
    .C(n_12595_o_0),
    .Y(n_12596_o_0));
 NAND2xp33_ASAP7_75t_R n_12597 (.A(key[36]),
    .B(ld),
    .Y(n_12597_o_0));
 OAI21xp33_ASAP7_75t_R n_12598 (.A1(ld),
    .A2(n_1885_o_0),
    .B(n_12597_o_0),
    .Y(n_12598_o_0));
 INVx1_ASAP7_75t_R n_12599 (.A(n_1876_o_0),
    .Y(n_12599_o_0));
 AOI21xp33_ASAP7_75t_R n_1260 (.A1(n_878_o_0),
    .A2(n_886_o_0),
    .B(n_1259_o_0),
    .Y(n_1260_o_0));
 NAND2xp33_ASAP7_75t_R n_12600 (.A(key[37]),
    .B(ld),
    .Y(n_12600_o_0));
 OAI21xp33_ASAP7_75t_R n_12601 (.A1(ld),
    .A2(n_12599_o_0),
    .B(n_12600_o_0),
    .Y(n_12601_o_0));
 INVx1_ASAP7_75t_R n_12602 (.A(n_1869_o_0),
    .Y(n_12602_o_0));
 NAND2xp33_ASAP7_75t_R n_12603 (.A(key[38]),
    .B(ld),
    .Y(n_12603_o_0));
 OAI21xp33_ASAP7_75t_R n_12604 (.A1(ld),
    .A2(n_12602_o_0),
    .B(n_12603_o_0),
    .Y(n_12604_o_0));
 INVx1_ASAP7_75t_R n_12605 (.A(n_1862_o_0),
    .Y(n_12605_o_0));
 NAND2xp33_ASAP7_75t_R n_12606 (.A(key[39]),
    .B(ld),
    .Y(n_12606_o_0));
 OAI21xp33_ASAP7_75t_R n_12607 (.A1(ld),
    .A2(n_12605_o_0),
    .B(n_12606_o_0),
    .Y(n_12607_o_0));
 XNOR2xp5_ASAP7_75t_R n_12608 (.A(_00932_),
    .B(n_1384_o_0),
    .Y(n_12608_o_0));
 NAND2xp33_ASAP7_75t_R n_12609 (.A(key[40]),
    .B(ld),
    .Y(n_12609_o_0));
 NAND3xp33_ASAP7_75t_R n_1261 (.A(n_1085_o_0),
    .B(n_944_o_0),
    .C(n_878_o_0),
    .Y(n_1261_o_0));
 OAI21xp33_ASAP7_75t_R n_12610 (.A1(ld),
    .A2(n_12608_o_0),
    .B(n_12609_o_0),
    .Y(n_12610_o_0));
 XNOR2xp5_ASAP7_75t_R n_12611 (.A(_00933_),
    .B(n_1375_o_0),
    .Y(n_12611_o_0));
 NAND2xp33_ASAP7_75t_R n_12612 (.A(key[41]),
    .B(ld),
    .Y(n_12612_o_0));
 OAI21xp33_ASAP7_75t_R n_12613 (.A1(ld),
    .A2(n_12611_o_0),
    .B(n_12612_o_0),
    .Y(n_12613_o_0));
 NAND2xp33_ASAP7_75t_R n_12614 (.A(ld),
    .B(text_in[0]),
    .Y(n_12614_o_0));
 OAI21xp33_ASAP7_75t_R n_12615 (.A1(_00411_),
    .A2(ld),
    .B(n_12614_o_0),
    .Y(n_12615_o_0));
 NAND2xp33_ASAP7_75t_R n_12616 (.A(ld),
    .B(text_in[1]),
    .Y(n_12616_o_0));
 OAI21xp33_ASAP7_75t_R n_12617 (.A1(_00410_),
    .A2(ld),
    .B(n_12616_o_0),
    .Y(n_12617_o_0));
 NAND2xp33_ASAP7_75t_R n_12618 (.A(ld),
    .B(text_in[2]),
    .Y(n_12618_o_0));
 OAI21xp33_ASAP7_75t_R n_12619 (.A1(_00413_),
    .A2(ld),
    .B(n_12618_o_0),
    .Y(n_12619_o_0));
 AOI21xp33_ASAP7_75t_R n_1262 (.A1(n_890_o_0),
    .A2(n_1261_o_0),
    .B(net16),
    .Y(n_1262_o_0));
 NAND2xp33_ASAP7_75t_R n_12620 (.A(ld),
    .B(text_in[3]),
    .Y(n_12620_o_0));
 OAI21xp33_ASAP7_75t_R n_12621 (.A1(_00728_),
    .A2(ld),
    .B(n_12620_o_0),
    .Y(n_12621_o_0));
 NAND2xp33_ASAP7_75t_R n_12622 (.A(ld),
    .B(text_in[4]),
    .Y(n_12622_o_0));
 OAI21xp33_ASAP7_75t_R n_12623 (.A1(_00727_),
    .A2(ld),
    .B(n_12622_o_0),
    .Y(n_12623_o_0));
 NAND2xp33_ASAP7_75t_R n_12624 (.A(ld),
    .B(text_in[5]),
    .Y(n_12624_o_0));
 OAI21xp33_ASAP7_75t_R n_12625 (.A1(_00726_),
    .A2(ld),
    .B(n_12624_o_0),
    .Y(n_12625_o_0));
 NAND2xp33_ASAP7_75t_R n_12626 (.A(ld),
    .B(text_in[6]),
    .Y(n_12626_o_0));
 OAI21xp33_ASAP7_75t_R n_12627 (.A1(_00725_),
    .A2(ld),
    .B(n_12626_o_0),
    .Y(n_12627_o_0));
 NAND2xp33_ASAP7_75t_R n_12628 (.A(ld),
    .B(text_in[7]),
    .Y(n_12628_o_0));
 OAI21xp33_ASAP7_75t_R n_12629 (.A1(_00724_),
    .A2(ld),
    .B(n_12628_o_0),
    .Y(n_12629_o_0));
 OAI21xp33_ASAP7_75t_R n_1263 (.A1(n_1260_o_0),
    .A2(n_1262_o_0),
    .B(n_903_o_0),
    .Y(n_1263_o_0));
 NAND2xp33_ASAP7_75t_R n_12630 (.A(ld),
    .B(text_in[8]),
    .Y(n_12630_o_0));
 OAI21xp33_ASAP7_75t_R n_12631 (.A1(_00606_),
    .A2(ld),
    .B(n_12630_o_0),
    .Y(n_12631_o_0));
 NAND2xp33_ASAP7_75t_R n_12632 (.A(ld),
    .B(text_in[9]),
    .Y(n_12632_o_0));
 OAI21xp33_ASAP7_75t_R n_12633 (.A1(_00605_),
    .A2(ld),
    .B(n_12632_o_0),
    .Y(n_12633_o_0));
 NAND2xp33_ASAP7_75t_R n_12634 (.A(ld),
    .B(text_in[10]),
    .Y(n_12634_o_0));
 OAI21xp33_ASAP7_75t_R n_12635 (.A1(_00608_),
    .A2(ld),
    .B(n_12634_o_0),
    .Y(n_12635_o_0));
 NAND2xp33_ASAP7_75t_R n_12636 (.A(ld),
    .B(text_in[11]),
    .Y(n_12636_o_0));
 OAI21xp33_ASAP7_75t_R n_12637 (.A1(_00723_),
    .A2(ld),
    .B(n_12636_o_0),
    .Y(n_12637_o_0));
 NAND2xp33_ASAP7_75t_R n_12638 (.A(ld),
    .B(text_in[12]),
    .Y(n_12638_o_0));
 OAI21xp33_ASAP7_75t_R n_12639 (.A1(_00722_),
    .A2(ld),
    .B(n_12638_o_0),
    .Y(n_12639_o_0));
 AOI21xp33_ASAP7_75t_R n_1264 (.A1(n_1258_o_0),
    .A2(n_1263_o_0),
    .B(n_972_o_0),
    .Y(n_1264_o_0));
 NAND2xp33_ASAP7_75t_R n_12640 (.A(ld),
    .B(text_in[13]),
    .Y(n_12640_o_0));
 OAI21xp33_ASAP7_75t_R n_12641 (.A1(_00721_),
    .A2(ld),
    .B(n_12640_o_0),
    .Y(n_12641_o_0));
 NAND2xp33_ASAP7_75t_R n_12642 (.A(ld),
    .B(text_in[14]),
    .Y(n_12642_o_0));
 OAI21xp33_ASAP7_75t_R n_12643 (.A1(_00720_),
    .A2(ld),
    .B(n_12642_o_0),
    .Y(n_12643_o_0));
 NAND2xp33_ASAP7_75t_R n_12644 (.A(ld),
    .B(text_in[15]),
    .Y(n_12644_o_0));
 OAI21xp33_ASAP7_75t_R n_12645 (.A1(_00719_),
    .A2(ld),
    .B(n_12644_o_0),
    .Y(n_12645_o_0));
 NAND2xp33_ASAP7_75t_R n_12646 (.A(ld),
    .B(text_in[16]),
    .Y(n_12646_o_0));
 OAI21xp33_ASAP7_75t_R n_12647 (.A1(_00560_),
    .A2(ld),
    .B(n_12646_o_0),
    .Y(n_12647_o_0));
 NAND2xp33_ASAP7_75t_R n_12648 (.A(ld),
    .B(text_in[17]),
    .Y(n_12648_o_0));
 OAI21xp33_ASAP7_75t_R n_12649 (.A1(_00559_),
    .A2(ld),
    .B(n_12648_o_0),
    .Y(n_12649_o_0));
 AOI31xp33_ASAP7_75t_R n_1265 (.A1(n_877_o_0),
    .A2(n_910_o_0),
    .A3(n_990_o_0),
    .B(net14),
    .Y(n_1265_o_0));
 NAND2xp33_ASAP7_75t_R n_12650 (.A(ld),
    .B(text_in[18]),
    .Y(n_12650_o_0));
 OAI21xp33_ASAP7_75t_R n_12651 (.A1(_00562_),
    .A2(ld),
    .B(n_12650_o_0),
    .Y(n_12651_o_0));
 NAND2xp33_ASAP7_75t_R n_12652 (.A(ld),
    .B(text_in[19]),
    .Y(n_12652_o_0));
 OAI21xp33_ASAP7_75t_R n_12653 (.A1(_00718_),
    .A2(ld),
    .B(n_12652_o_0),
    .Y(n_12653_o_0));
 NAND2xp33_ASAP7_75t_R n_12654 (.A(ld),
    .B(text_in[20]),
    .Y(n_12654_o_0));
 OAI21xp33_ASAP7_75t_R n_12655 (.A1(_00717_),
    .A2(ld),
    .B(n_12654_o_0),
    .Y(n_12655_o_0));
 NAND2xp33_ASAP7_75t_R n_12656 (.A(ld),
    .B(text_in[21]),
    .Y(n_12656_o_0));
 OAI21xp33_ASAP7_75t_R n_12657 (.A1(_00716_),
    .A2(ld),
    .B(n_12656_o_0),
    .Y(n_12657_o_0));
 NAND2xp33_ASAP7_75t_R n_12658 (.A(ld),
    .B(text_in[22]),
    .Y(n_12658_o_0));
 OAI21xp33_ASAP7_75t_R n_12659 (.A1(_00715_),
    .A2(ld),
    .B(n_12658_o_0),
    .Y(n_12659_o_0));
 OAI21xp33_ASAP7_75t_R n_1266 (.A1(n_1006_o_0),
    .A2(n_1167_o_0),
    .B(n_891_o_0),
    .Y(n_1266_o_0));
 NAND2xp33_ASAP7_75t_R n_12660 (.A(ld),
    .B(text_in[23]),
    .Y(n_12660_o_0));
 OAI21xp33_ASAP7_75t_R n_12661 (.A1(_00714_),
    .A2(ld),
    .B(n_12660_o_0),
    .Y(n_12661_o_0));
 NAND2xp33_ASAP7_75t_R n_12662 (.A(ld),
    .B(text_in[24]),
    .Y(n_12662_o_0));
 OAI21xp33_ASAP7_75t_R n_12663 (.A1(_00520_),
    .A2(ld),
    .B(n_12662_o_0),
    .Y(n_12663_o_0));
 NAND2xp33_ASAP7_75t_R n_12664 (.A(ld),
    .B(text_in[25]),
    .Y(n_12664_o_0));
 OAI21xp33_ASAP7_75t_R n_12665 (.A1(_00519_),
    .A2(ld),
    .B(n_12664_o_0),
    .Y(n_12665_o_0));
 NAND2xp33_ASAP7_75t_R n_12666 (.A(ld),
    .B(text_in[26]),
    .Y(n_12666_o_0));
 OAI21xp33_ASAP7_75t_R n_12667 (.A1(_00522_),
    .A2(ld),
    .B(n_12666_o_0),
    .Y(n_12667_o_0));
 NAND2xp33_ASAP7_75t_R n_12668 (.A(ld),
    .B(text_in[27]),
    .Y(n_12668_o_0));
 OAI21xp33_ASAP7_75t_R n_12669 (.A1(_00713_),
    .A2(ld),
    .B(n_12668_o_0),
    .Y(n_12669_o_0));
 NOR3xp33_ASAP7_75t_R n_1267 (.A(n_913_o_0),
    .B(n_877_o_0),
    .C(n_881_o_0),
    .Y(n_1267_o_0));
 NAND2xp33_ASAP7_75t_R n_12670 (.A(ld),
    .B(text_in[28]),
    .Y(n_12670_o_0));
 OAI21xp33_ASAP7_75t_R n_12671 (.A1(_00712_),
    .A2(ld),
    .B(n_12670_o_0),
    .Y(n_12671_o_0));
 NAND2xp33_ASAP7_75t_R n_12672 (.A(ld),
    .B(text_in[29]),
    .Y(n_12672_o_0));
 OAI21xp33_ASAP7_75t_R n_12673 (.A1(_00711_),
    .A2(ld),
    .B(n_12672_o_0),
    .Y(n_12673_o_0));
 NAND2xp33_ASAP7_75t_R n_12674 (.A(ld),
    .B(text_in[30]),
    .Y(n_12674_o_0));
 OAI21xp33_ASAP7_75t_R n_12675 (.A1(_00710_),
    .A2(ld),
    .B(n_12674_o_0),
    .Y(n_12675_o_0));
 NAND2xp33_ASAP7_75t_R n_12676 (.A(ld),
    .B(text_in[31]),
    .Y(n_12676_o_0));
 OAI21xp33_ASAP7_75t_R n_12677 (.A1(_00709_),
    .A2(ld),
    .B(n_12676_o_0),
    .Y(n_12677_o_0));
 NAND2xp33_ASAP7_75t_R n_12678 (.A(ld),
    .B(text_in[32]),
    .Y(n_12678_o_0));
 OAI21xp33_ASAP7_75t_R n_12679 (.A1(_00638_),
    .A2(ld),
    .B(n_12678_o_0),
    .Y(n_12679_o_0));
 OAI31xp33_ASAP7_75t_R n_1268 (.A1(n_1150_o_0),
    .A2(n_1266_o_0),
    .A3(n_1267_o_0),
    .B(n_903_o_0),
    .Y(n_1268_o_0));
 NAND2xp33_ASAP7_75t_R n_12680 (.A(ld),
    .B(text_in[33]),
    .Y(n_12680_o_0));
 OAI21xp33_ASAP7_75t_R n_12681 (.A1(_00637_),
    .A2(ld),
    .B(n_12680_o_0),
    .Y(n_12681_o_0));
 NAND2xp33_ASAP7_75t_R n_12682 (.A(ld),
    .B(text_in[34]),
    .Y(n_12682_o_0));
 OAI21xp33_ASAP7_75t_R n_12683 (.A1(_00639_),
    .A2(ld),
    .B(n_12682_o_0),
    .Y(n_12683_o_0));
 NAND2xp33_ASAP7_75t_R n_12684 (.A(ld),
    .B(text_in[35]),
    .Y(n_12684_o_0));
 OAI21xp33_ASAP7_75t_R n_12685 (.A1(_00708_),
    .A2(ld),
    .B(n_12684_o_0),
    .Y(n_12685_o_0));
 NAND2xp33_ASAP7_75t_R n_12686 (.A(ld),
    .B(text_in[36]),
    .Y(n_12686_o_0));
 OAI21xp33_ASAP7_75t_R n_12687 (.A1(_00707_),
    .A2(ld),
    .B(n_12686_o_0),
    .Y(n_12687_o_0));
 NAND2xp33_ASAP7_75t_R n_12688 (.A(ld),
    .B(text_in[37]),
    .Y(n_12688_o_0));
 OAI21xp33_ASAP7_75t_R n_12689 (.A1(_00706_),
    .A2(ld),
    .B(n_12688_o_0),
    .Y(n_12689_o_0));
 AOI21xp33_ASAP7_75t_R n_1269 (.A1(n_1156_o_0),
    .A2(n_1265_o_0),
    .B(n_1268_o_0),
    .Y(n_1269_o_0));
 NAND2xp33_ASAP7_75t_R n_12690 (.A(ld),
    .B(text_in[38]),
    .Y(n_12690_o_0));
 OAI21xp33_ASAP7_75t_R n_12691 (.A1(_00705_),
    .A2(ld),
    .B(n_12690_o_0),
    .Y(n_12691_o_0));
 NAND2xp33_ASAP7_75t_R n_12692 (.A(ld),
    .B(text_in[39]),
    .Y(n_12692_o_0));
 OAI21xp33_ASAP7_75t_R n_12693 (.A1(_00704_),
    .A2(ld),
    .B(n_12692_o_0),
    .Y(n_12693_o_0));
 NAND2xp33_ASAP7_75t_R n_12694 (.A(ld),
    .B(text_in[40]),
    .Y(n_12694_o_0));
 OAI21xp33_ASAP7_75t_R n_12695 (.A1(_00594_),
    .A2(ld),
    .B(n_12694_o_0),
    .Y(n_12695_o_0));
 NAND2xp33_ASAP7_75t_R n_12696 (.A(ld),
    .B(text_in[41]),
    .Y(n_12696_o_0));
 OAI21xp33_ASAP7_75t_R n_12697 (.A1(_00593_),
    .A2(ld),
    .B(n_12696_o_0),
    .Y(n_12697_o_0));
 NAND2xp33_ASAP7_75t_R n_12698 (.A(ld),
    .B(text_in[42]),
    .Y(n_12698_o_0));
 OAI21xp33_ASAP7_75t_R n_12699 (.A1(_00596_),
    .A2(ld),
    .B(n_12698_o_0),
    .Y(n_12699_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1270 (.A1(n_860_o_0),
    .A2(net32),
    .B(n_982_o_0),
    .C(n_878_o_0),
    .Y(n_1270_o_0));
 NAND2xp33_ASAP7_75t_R n_12700 (.A(ld),
    .B(text_in[43]),
    .Y(n_12700_o_0));
 OAI21xp33_ASAP7_75t_R n_12701 (.A1(_00703_),
    .A2(ld),
    .B(n_12700_o_0),
    .Y(n_12701_o_0));
 NAND2xp33_ASAP7_75t_R n_12702 (.A(ld),
    .B(text_in[44]),
    .Y(n_12702_o_0));
 OAI21xp33_ASAP7_75t_R n_12703 (.A1(_00702_),
    .A2(ld),
    .B(n_12702_o_0),
    .Y(n_12703_o_0));
 NAND2xp33_ASAP7_75t_R n_12704 (.A(ld),
    .B(text_in[45]),
    .Y(n_12704_o_0));
 OAI21xp33_ASAP7_75t_R n_12705 (.A1(_00701_),
    .A2(ld),
    .B(n_12704_o_0),
    .Y(n_12705_o_0));
 NAND2xp33_ASAP7_75t_R n_12706 (.A(ld),
    .B(text_in[46]),
    .Y(n_12706_o_0));
 OAI21xp33_ASAP7_75t_R n_12707 (.A1(_00700_),
    .A2(ld),
    .B(n_12706_o_0),
    .Y(n_12707_o_0));
 NAND2xp33_ASAP7_75t_R n_12708 (.A(ld),
    .B(text_in[47]),
    .Y(n_12708_o_0));
 OAI21xp33_ASAP7_75t_R n_12709 (.A1(_00699_),
    .A2(ld),
    .B(n_12708_o_0),
    .Y(n_12709_o_0));
 OAI21xp33_ASAP7_75t_R n_1271 (.A1(n_847_o_0),
    .A2(n_877_o_0),
    .B(n_864_o_0),
    .Y(n_1271_o_0));
 NAND2xp33_ASAP7_75t_R n_12710 (.A(ld),
    .B(text_in[48]),
    .Y(n_12710_o_0));
 OAI21xp33_ASAP7_75t_R n_12711 (.A1(_00550_),
    .A2(ld),
    .B(n_12710_o_0),
    .Y(n_12711_o_0));
 NAND2xp33_ASAP7_75t_R n_12712 (.A(ld),
    .B(text_in[49]),
    .Y(n_12712_o_0));
 OAI21xp33_ASAP7_75t_R n_12713 (.A1(_00549_),
    .A2(ld),
    .B(n_12712_o_0),
    .Y(n_12713_o_0));
 NAND2xp33_ASAP7_75t_R n_12714 (.A(ld),
    .B(text_in[50]),
    .Y(n_12714_o_0));
 OAI21xp33_ASAP7_75t_R n_12715 (.A1(_00552_),
    .A2(ld),
    .B(n_12714_o_0),
    .Y(n_12715_o_0));
 NAND2xp33_ASAP7_75t_R n_12716 (.A(ld),
    .B(text_in[51]),
    .Y(n_12716_o_0));
 OAI21xp33_ASAP7_75t_R n_12717 (.A1(_00698_),
    .A2(ld),
    .B(n_12716_o_0),
    .Y(n_12717_o_0));
 NAND2xp33_ASAP7_75t_R n_12718 (.A(ld),
    .B(text_in[52]),
    .Y(n_12718_o_0));
 OAI21xp33_ASAP7_75t_R n_12719 (.A1(_00697_),
    .A2(ld),
    .B(n_12718_o_0),
    .Y(n_12719_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1272 (.A1(n_877_o_0),
    .A2(n_956_o_0),
    .B(n_1271_o_0),
    .C(net42),
    .Y(n_1272_o_0));
 NAND2xp33_ASAP7_75t_R n_12720 (.A(ld),
    .B(text_in[53]),
    .Y(n_12720_o_0));
 OAI21xp33_ASAP7_75t_R n_12721 (.A1(_00696_),
    .A2(ld),
    .B(n_12720_o_0),
    .Y(n_12721_o_0));
 NAND2xp33_ASAP7_75t_R n_12722 (.A(ld),
    .B(text_in[54]),
    .Y(n_12722_o_0));
 OAI21xp33_ASAP7_75t_R n_12723 (.A1(_00695_),
    .A2(ld),
    .B(n_12722_o_0),
    .Y(n_12723_o_0));
 NAND2xp33_ASAP7_75t_R n_12724 (.A(ld),
    .B(text_in[55]),
    .Y(n_12724_o_0));
 OAI21xp33_ASAP7_75t_R n_12725 (.A1(_00694_),
    .A2(ld),
    .B(n_12724_o_0),
    .Y(n_12725_o_0));
 NAND2xp33_ASAP7_75t_R n_12726 (.A(ld),
    .B(text_in[56]),
    .Y(n_12726_o_0));
 OAI21xp33_ASAP7_75t_R n_12727 (.A1(_00510_),
    .A2(ld),
    .B(n_12726_o_0),
    .Y(n_12727_o_0));
 NAND2xp33_ASAP7_75t_R n_12728 (.A(ld),
    .B(text_in[57]),
    .Y(n_12728_o_0));
 OAI21xp33_ASAP7_75t_R n_12729 (.A1(_00509_),
    .A2(ld),
    .B(n_12728_o_0),
    .Y(n_12729_o_0));
 AOI311xp33_ASAP7_75t_R n_1273 (.A1(net16),
    .A2(n_1189_o_0),
    .A3(n_1270_o_0),
    .B(n_903_o_0),
    .C(n_1272_o_0),
    .Y(n_1273_o_0));
 NAND2xp33_ASAP7_75t_R n_12730 (.A(ld),
    .B(text_in[58]),
    .Y(n_12730_o_0));
 OAI21xp33_ASAP7_75t_R n_12731 (.A1(_00512_),
    .A2(ld),
    .B(n_12730_o_0),
    .Y(n_12731_o_0));
 NAND2xp33_ASAP7_75t_R n_12732 (.A(ld),
    .B(text_in[59]),
    .Y(n_12732_o_0));
 OAI21xp33_ASAP7_75t_R n_12733 (.A1(_00693_),
    .A2(ld),
    .B(n_12732_o_0),
    .Y(n_12733_o_0));
 NAND2xp33_ASAP7_75t_R n_12734 (.A(ld),
    .B(text_in[60]),
    .Y(n_12734_o_0));
 OAI21xp33_ASAP7_75t_R n_12735 (.A1(_00692_),
    .A2(ld),
    .B(n_12734_o_0),
    .Y(n_12735_o_0));
 NAND2xp33_ASAP7_75t_R n_12736 (.A(ld),
    .B(text_in[61]),
    .Y(n_12736_o_0));
 OAI21xp33_ASAP7_75t_R n_12737 (.A1(_00691_),
    .A2(ld),
    .B(n_12736_o_0),
    .Y(n_12737_o_0));
 NAND2xp33_ASAP7_75t_R n_12738 (.A(ld),
    .B(text_in[62]),
    .Y(n_12738_o_0));
 OAI21xp33_ASAP7_75t_R n_12739 (.A1(_00690_),
    .A2(ld),
    .B(n_12738_o_0),
    .Y(n_12739_o_0));
 NOR3xp33_ASAP7_75t_R n_1274 (.A(n_1269_o_0),
    .B(n_971_o_0),
    .C(n_1273_o_0),
    .Y(n_1274_o_0));
 NAND2xp33_ASAP7_75t_R n_12740 (.A(ld),
    .B(text_in[63]),
    .Y(n_12740_o_0));
 OAI21xp33_ASAP7_75t_R n_12741 (.A1(_00689_),
    .A2(ld),
    .B(n_12740_o_0),
    .Y(n_12741_o_0));
 NAND2xp33_ASAP7_75t_R n_12742 (.A(ld),
    .B(text_in[64]),
    .Y(n_12742_o_0));
 OAI21xp33_ASAP7_75t_R n_12743 (.A1(_00628_),
    .A2(ld),
    .B(n_12742_o_0),
    .Y(n_12743_o_0));
 NAND2xp33_ASAP7_75t_R n_12744 (.A(ld),
    .B(text_in[65]),
    .Y(n_12744_o_0));
 OAI21xp33_ASAP7_75t_R n_12745 (.A1(_00627_),
    .A2(ld),
    .B(n_12744_o_0),
    .Y(n_12745_o_0));
 NAND2xp33_ASAP7_75t_R n_12746 (.A(ld),
    .B(text_in[66]),
    .Y(n_12746_o_0));
 OAI21xp33_ASAP7_75t_R n_12747 (.A1(_00630_),
    .A2(ld),
    .B(n_12746_o_0),
    .Y(n_12747_o_0));
 NAND2xp33_ASAP7_75t_R n_12748 (.A(ld),
    .B(text_in[67]),
    .Y(n_12748_o_0));
 OAI21xp33_ASAP7_75t_R n_12749 (.A1(_00688_),
    .A2(ld),
    .B(n_12748_o_0),
    .Y(n_12749_o_0));
 OAI21xp33_ASAP7_75t_R n_1275 (.A1(n_915_o_0),
    .A2(n_890_o_0),
    .B(n_891_o_0),
    .Y(n_1275_o_0));
 NAND2xp33_ASAP7_75t_R n_12750 (.A(ld),
    .B(text_in[68]),
    .Y(n_12750_o_0));
 OAI21xp33_ASAP7_75t_R n_12751 (.A1(_00687_),
    .A2(ld),
    .B(n_12750_o_0),
    .Y(n_12751_o_0));
 NAND2xp33_ASAP7_75t_R n_12752 (.A(ld),
    .B(text_in[69]),
    .Y(n_12752_o_0));
 OAI21xp33_ASAP7_75t_R n_12753 (.A1(_00686_),
    .A2(ld),
    .B(n_12752_o_0),
    .Y(n_12753_o_0));
 NAND2xp33_ASAP7_75t_R n_12754 (.A(ld),
    .B(text_in[70]),
    .Y(n_12754_o_0));
 OAI21xp33_ASAP7_75t_R n_12755 (.A1(_00685_),
    .A2(ld),
    .B(n_12754_o_0),
    .Y(n_12755_o_0));
 NAND2xp33_ASAP7_75t_R n_12756 (.A(ld),
    .B(text_in[71]),
    .Y(n_12756_o_0));
 OAI21xp33_ASAP7_75t_R n_12757 (.A1(_00684_),
    .A2(ld),
    .B(n_12756_o_0),
    .Y(n_12757_o_0));
 NAND2xp33_ASAP7_75t_R n_12758 (.A(ld),
    .B(text_in[72]),
    .Y(n_12758_o_0));
 OAI21xp33_ASAP7_75t_R n_12759 (.A1(_00582_),
    .A2(ld),
    .B(n_12758_o_0),
    .Y(n_12759_o_0));
 AOI21xp33_ASAP7_75t_R n_1276 (.A1(n_882_o_0),
    .A2(n_954_o_0),
    .B(n_891_o_0),
    .Y(n_1276_o_0));
 NAND2xp33_ASAP7_75t_R n_12760 (.A(ld),
    .B(text_in[73]),
    .Y(n_12760_o_0));
 OAI21xp33_ASAP7_75t_R n_12761 (.A1(_00581_),
    .A2(ld),
    .B(n_12760_o_0),
    .Y(n_12761_o_0));
 NAND2xp33_ASAP7_75t_R n_12762 (.A(ld),
    .B(text_in[74]),
    .Y(n_12762_o_0));
 OAI21xp33_ASAP7_75t_R n_12763 (.A1(_00584_),
    .A2(ld),
    .B(n_12762_o_0),
    .Y(n_12763_o_0));
 NAND2xp33_ASAP7_75t_R n_12764 (.A(ld),
    .B(text_in[75]),
    .Y(n_12764_o_0));
 OAI21xp33_ASAP7_75t_R n_12765 (.A1(_00683_),
    .A2(ld),
    .B(n_12764_o_0),
    .Y(n_12765_o_0));
 NAND2xp33_ASAP7_75t_R n_12766 (.A(ld),
    .B(text_in[76]),
    .Y(n_12766_o_0));
 OAI21xp33_ASAP7_75t_R n_12767 (.A1(_00682_),
    .A2(ld),
    .B(n_12766_o_0),
    .Y(n_12767_o_0));
 NAND2xp33_ASAP7_75t_R n_12768 (.A(ld),
    .B(text_in[77]),
    .Y(n_12768_o_0));
 OAI21xp33_ASAP7_75t_R n_12769 (.A1(_00681_),
    .A2(ld),
    .B(n_12768_o_0),
    .Y(n_12769_o_0));
 OAI21xp33_ASAP7_75t_R n_1277 (.A1(n_877_o_0),
    .A2(n_989_o_0),
    .B(n_1276_o_0),
    .Y(n_1277_o_0));
 NAND2xp33_ASAP7_75t_R n_12770 (.A(ld),
    .B(text_in[78]),
    .Y(n_12770_o_0));
 OAI21xp33_ASAP7_75t_R n_12771 (.A1(_00680_),
    .A2(ld),
    .B(n_12770_o_0),
    .Y(n_12771_o_0));
 NAND2xp33_ASAP7_75t_R n_12772 (.A(ld),
    .B(text_in[79]),
    .Y(n_12772_o_0));
 OAI21xp33_ASAP7_75t_R n_12773 (.A1(_00679_),
    .A2(ld),
    .B(n_12772_o_0),
    .Y(n_12773_o_0));
 NAND2xp33_ASAP7_75t_R n_12774 (.A(ld),
    .B(text_in[80]),
    .Y(n_12774_o_0));
 OAI21xp33_ASAP7_75t_R n_12775 (.A1(_00540_),
    .A2(ld),
    .B(n_12774_o_0),
    .Y(n_12775_o_0));
 NAND2xp33_ASAP7_75t_R n_12776 (.A(ld),
    .B(text_in[81]),
    .Y(n_12776_o_0));
 OAI21xp33_ASAP7_75t_R n_12777 (.A1(_00539_),
    .A2(ld),
    .B(n_12776_o_0),
    .Y(n_12777_o_0));
 NAND2xp33_ASAP7_75t_R n_12778 (.A(ld),
    .B(text_in[82]),
    .Y(n_12778_o_0));
 OAI21xp33_ASAP7_75t_R n_12779 (.A1(_00542_),
    .A2(ld),
    .B(n_12778_o_0),
    .Y(n_12779_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1278 (.A1(n_943_o_0),
    .A2(n_953_o_0),
    .B(n_1275_o_0),
    .C(n_1277_o_0),
    .Y(n_1278_o_0));
 NAND2xp33_ASAP7_75t_R n_12780 (.A(ld),
    .B(text_in[83]),
    .Y(n_12780_o_0));
 OAI21xp33_ASAP7_75t_R n_12781 (.A1(_00678_),
    .A2(ld),
    .B(n_12780_o_0),
    .Y(n_12781_o_0));
 NAND2xp33_ASAP7_75t_R n_12782 (.A(ld),
    .B(text_in[84]),
    .Y(n_12782_o_0));
 OAI21xp33_ASAP7_75t_R n_12783 (.A1(_00677_),
    .A2(ld),
    .B(n_12782_o_0),
    .Y(n_12783_o_0));
 NAND2xp33_ASAP7_75t_R n_12784 (.A(ld),
    .B(text_in[85]),
    .Y(n_12784_o_0));
 OAI21xp33_ASAP7_75t_R n_12785 (.A1(_00676_),
    .A2(ld),
    .B(n_12784_o_0),
    .Y(n_12785_o_0));
 NAND2xp33_ASAP7_75t_R n_12786 (.A(ld),
    .B(text_in[86]),
    .Y(n_12786_o_0));
 OAI21xp33_ASAP7_75t_R n_12787 (.A1(_00675_),
    .A2(ld),
    .B(n_12786_o_0),
    .Y(n_12787_o_0));
 NAND2xp33_ASAP7_75t_R n_12788 (.A(ld),
    .B(text_in[87]),
    .Y(n_12788_o_0));
 OAI21xp33_ASAP7_75t_R n_12789 (.A1(_00674_),
    .A2(ld),
    .B(n_12788_o_0),
    .Y(n_12789_o_0));
 OAI21xp33_ASAP7_75t_R n_1279 (.A1(n_887_o_0),
    .A2(n_1004_o_0),
    .B(net42),
    .Y(n_1279_o_0));
 NAND2xp33_ASAP7_75t_R n_12790 (.A(ld),
    .B(text_in[88]),
    .Y(n_12790_o_0));
 OAI21xp33_ASAP7_75t_R n_12791 (.A1(_00500_),
    .A2(ld),
    .B(n_12790_o_0),
    .Y(n_12791_o_0));
 NAND2xp33_ASAP7_75t_R n_12792 (.A(ld),
    .B(text_in[89]),
    .Y(n_12792_o_0));
 OAI21xp33_ASAP7_75t_R n_12793 (.A1(_00499_),
    .A2(ld),
    .B(n_12792_o_0),
    .Y(n_12793_o_0));
 NAND2xp33_ASAP7_75t_R n_12794 (.A(ld),
    .B(text_in[90]),
    .Y(n_12794_o_0));
 OAI21xp33_ASAP7_75t_R n_12795 (.A1(_00502_),
    .A2(ld),
    .B(n_12794_o_0),
    .Y(n_12795_o_0));
 NAND2xp33_ASAP7_75t_R n_12796 (.A(ld),
    .B(text_in[91]),
    .Y(n_12796_o_0));
 OAI21xp33_ASAP7_75t_R n_12797 (.A1(_00673_),
    .A2(ld),
    .B(n_12796_o_0),
    .Y(n_12797_o_0));
 NAND2xp33_ASAP7_75t_R n_12798 (.A(ld),
    .B(text_in[92]),
    .Y(n_12798_o_0));
 OAI21xp33_ASAP7_75t_R n_12799 (.A1(_00672_),
    .A2(ld),
    .B(n_12798_o_0),
    .Y(n_12799_o_0));
 AOI31xp33_ASAP7_75t_R n_1280 (.A1(n_877_o_0),
    .A2(n_990_o_0),
    .A3(n_910_o_0),
    .B(n_829_o_0),
    .Y(n_1280_o_0));
 NAND2xp33_ASAP7_75t_R n_12800 (.A(ld),
    .B(text_in[93]),
    .Y(n_12800_o_0));
 OAI21xp33_ASAP7_75t_R n_12801 (.A1(_00671_),
    .A2(ld),
    .B(n_12800_o_0),
    .Y(n_12801_o_0));
 NAND2xp33_ASAP7_75t_R n_12802 (.A(ld),
    .B(text_in[94]),
    .Y(n_12802_o_0));
 OAI21xp33_ASAP7_75t_R n_12803 (.A1(_00670_),
    .A2(ld),
    .B(n_12802_o_0),
    .Y(n_12803_o_0));
 NAND2xp33_ASAP7_75t_R n_12804 (.A(ld),
    .B(text_in[95]),
    .Y(n_12804_o_0));
 OAI21xp33_ASAP7_75t_R n_12805 (.A1(_00669_),
    .A2(ld),
    .B(n_12804_o_0),
    .Y(n_12805_o_0));
 NAND2xp33_ASAP7_75t_R n_12806 (.A(ld),
    .B(text_in[96]),
    .Y(n_12806_o_0));
 OAI21xp33_ASAP7_75t_R n_12807 (.A1(_00618_),
    .A2(ld),
    .B(n_12806_o_0),
    .Y(n_12807_o_0));
 NAND2xp33_ASAP7_75t_R n_12808 (.A(ld),
    .B(text_in[97]),
    .Y(n_12808_o_0));
 OAI21xp33_ASAP7_75t_R n_12809 (.A1(_00617_),
    .A2(ld),
    .B(n_12808_o_0),
    .Y(n_12809_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1281 (.A1(n_1004_o_0),
    .A2(n_994_o_0),
    .B(n_1280_o_0),
    .C(n_904_o_0),
    .Y(n_1281_o_0));
 NAND2xp33_ASAP7_75t_R n_12810 (.A(ld),
    .B(text_in[98]),
    .Y(n_12810_o_0));
 OAI21xp33_ASAP7_75t_R n_12811 (.A1(_00620_),
    .A2(ld),
    .B(n_12810_o_0),
    .Y(n_12811_o_0));
 NAND2xp33_ASAP7_75t_R n_12812 (.A(ld),
    .B(text_in[99]),
    .Y(n_12812_o_0));
 OAI21xp33_ASAP7_75t_R n_12813 (.A1(_00668_),
    .A2(ld),
    .B(n_12812_o_0),
    .Y(n_12813_o_0));
 NAND2xp33_ASAP7_75t_R n_12814 (.A(ld),
    .B(text_in[100]),
    .Y(n_12814_o_0));
 OAI21xp33_ASAP7_75t_R n_12815 (.A1(_00667_),
    .A2(ld),
    .B(n_12814_o_0),
    .Y(n_12815_o_0));
 NAND2xp33_ASAP7_75t_R n_12816 (.A(ld),
    .B(text_in[101]),
    .Y(n_12816_o_0));
 OAI21xp33_ASAP7_75t_R n_12817 (.A1(_00666_),
    .A2(ld),
    .B(n_12816_o_0),
    .Y(n_12817_o_0));
 NAND2xp33_ASAP7_75t_R n_12818 (.A(ld),
    .B(text_in[102]),
    .Y(n_12818_o_0));
 OAI21xp33_ASAP7_75t_R n_12819 (.A1(_00665_),
    .A2(ld),
    .B(n_12818_o_0),
    .Y(n_12819_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1282 (.A1(n_866_o_0),
    .A2(n_877_o_0),
    .B(n_1279_o_0),
    .C(n_1281_o_0),
    .Y(n_1282_o_0));
 NAND2xp33_ASAP7_75t_R n_12820 (.A(ld),
    .B(text_in[103]),
    .Y(n_12820_o_0));
 OAI21xp33_ASAP7_75t_R n_12821 (.A1(_00664_),
    .A2(ld),
    .B(n_12820_o_0),
    .Y(n_12821_o_0));
 NAND2xp33_ASAP7_75t_R n_12822 (.A(ld),
    .B(text_in[104]),
    .Y(n_12822_o_0));
 OAI21xp33_ASAP7_75t_R n_12823 (.A1(_00570_),
    .A2(ld),
    .B(n_12822_o_0),
    .Y(n_12823_o_0));
 NAND2xp33_ASAP7_75t_R n_12824 (.A(ld),
    .B(text_in[105]),
    .Y(n_12824_o_0));
 OAI21xp33_ASAP7_75t_R n_12825 (.A1(_00569_),
    .A2(ld),
    .B(n_12824_o_0),
    .Y(n_12825_o_0));
 NAND2xp33_ASAP7_75t_R n_12826 (.A(ld),
    .B(text_in[106]),
    .Y(n_12826_o_0));
 OAI21xp33_ASAP7_75t_R n_12827 (.A1(_00572_),
    .A2(ld),
    .B(n_12826_o_0),
    .Y(n_12827_o_0));
 NAND2xp33_ASAP7_75t_R n_12828 (.A(ld),
    .B(text_in[107]),
    .Y(n_12828_o_0));
 OAI21xp33_ASAP7_75t_R n_12829 (.A1(_00663_),
    .A2(ld),
    .B(n_12828_o_0),
    .Y(n_12829_o_0));
 OAI21xp33_ASAP7_75t_R n_1283 (.A1(n_903_o_0),
    .A2(n_1278_o_0),
    .B(n_1282_o_0),
    .Y(n_1283_o_0));
 NAND2xp33_ASAP7_75t_R n_12830 (.A(ld),
    .B(text_in[108]),
    .Y(n_12830_o_0));
 OAI21xp33_ASAP7_75t_R n_12831 (.A1(_00662_),
    .A2(ld),
    .B(n_12830_o_0),
    .Y(n_12831_o_0));
 NAND2xp33_ASAP7_75t_R n_12832 (.A(ld),
    .B(text_in[109]),
    .Y(n_12832_o_0));
 OAI21xp33_ASAP7_75t_R n_12833 (.A1(_00661_),
    .A2(ld),
    .B(n_12832_o_0),
    .Y(n_12833_o_0));
 NAND2xp33_ASAP7_75t_R n_12834 (.A(ld),
    .B(text_in[110]),
    .Y(n_12834_o_0));
 OAI21xp33_ASAP7_75t_R n_12835 (.A1(_00660_),
    .A2(ld),
    .B(n_12834_o_0),
    .Y(n_12835_o_0));
 NAND2xp33_ASAP7_75t_R n_12836 (.A(ld),
    .B(text_in[111]),
    .Y(n_12836_o_0));
 OAI21xp33_ASAP7_75t_R n_12837 (.A1(_00659_),
    .A2(ld),
    .B(n_12836_o_0),
    .Y(n_12837_o_0));
 NAND2xp33_ASAP7_75t_R n_12838 (.A(ld),
    .B(text_in[112]),
    .Y(n_12838_o_0));
 OAI21xp33_ASAP7_75t_R n_12839 (.A1(_00530_),
    .A2(ld),
    .B(n_12838_o_0),
    .Y(n_12839_o_0));
 INVx1_ASAP7_75t_R n_1284 (.A(n_1074_o_0),
    .Y(n_1284_o_0));
 NAND2xp33_ASAP7_75t_R n_12840 (.A(ld),
    .B(text_in[113]),
    .Y(n_12840_o_0));
 OAI21xp33_ASAP7_75t_R n_12841 (.A1(_00529_),
    .A2(ld),
    .B(n_12840_o_0),
    .Y(n_12841_o_0));
 NAND2xp33_ASAP7_75t_R n_12842 (.A(ld),
    .B(text_in[114]),
    .Y(n_12842_o_0));
 OAI21xp33_ASAP7_75t_R n_12843 (.A1(_00532_),
    .A2(ld),
    .B(n_12842_o_0),
    .Y(n_12843_o_0));
 NAND2xp33_ASAP7_75t_R n_12844 (.A(ld),
    .B(text_in[115]),
    .Y(n_12844_o_0));
 OAI21xp33_ASAP7_75t_R n_12845 (.A1(_00658_),
    .A2(ld),
    .B(n_12844_o_0),
    .Y(n_12845_o_0));
 NAND2xp33_ASAP7_75t_R n_12846 (.A(ld),
    .B(text_in[116]),
    .Y(n_12846_o_0));
 OAI21xp33_ASAP7_75t_R n_12847 (.A1(_00657_),
    .A2(ld),
    .B(n_12846_o_0),
    .Y(n_12847_o_0));
 NAND2xp33_ASAP7_75t_R n_12848 (.A(ld),
    .B(text_in[117]),
    .Y(n_12848_o_0));
 OAI21xp33_ASAP7_75t_R n_12849 (.A1(_00656_),
    .A2(ld),
    .B(n_12848_o_0),
    .Y(n_12849_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1285 (.A1(n_1284_o_0),
    .A2(n_878_o_0),
    .B(net16),
    .C(n_903_o_0),
    .Y(n_1285_o_0));
 NAND2xp33_ASAP7_75t_R n_12850 (.A(ld),
    .B(text_in[118]),
    .Y(n_12850_o_0));
 OAI21xp33_ASAP7_75t_R n_12851 (.A1(_00655_),
    .A2(ld),
    .B(n_12850_o_0),
    .Y(n_12851_o_0));
 NAND2xp33_ASAP7_75t_R n_12852 (.A(ld),
    .B(text_in[119]),
    .Y(n_12852_o_0));
 OAI21xp33_ASAP7_75t_R n_12853 (.A1(_00654_),
    .A2(ld),
    .B(n_12852_o_0),
    .Y(n_12853_o_0));
 NAND2xp33_ASAP7_75t_R n_12854 (.A(ld),
    .B(text_in[120]),
    .Y(n_12854_o_0));
 OAI21xp33_ASAP7_75t_R n_12855 (.A1(_00490_),
    .A2(ld),
    .B(n_12854_o_0),
    .Y(n_12855_o_0));
 NAND2xp33_ASAP7_75t_R n_12856 (.A(ld),
    .B(text_in[121]),
    .Y(n_12856_o_0));
 OAI21xp33_ASAP7_75t_R n_12857 (.A1(_00489_),
    .A2(ld),
    .B(n_12856_o_0),
    .Y(n_12857_o_0));
 NAND2xp33_ASAP7_75t_R n_12858 (.A(ld),
    .B(text_in[122]),
    .Y(n_12858_o_0));
 OAI21xp33_ASAP7_75t_R n_12859 (.A1(_00492_),
    .A2(ld),
    .B(n_12858_o_0),
    .Y(n_12859_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1286 (.A1(n_878_o_0),
    .A2(n_1146_o_0),
    .B(n_1200_o_0),
    .C(n_891_o_0),
    .Y(n_1286_o_0));
 NAND2xp33_ASAP7_75t_R n_12860 (.A(ld),
    .B(text_in[123]),
    .Y(n_12860_o_0));
 OAI21xp33_ASAP7_75t_R n_12861 (.A1(_00653_),
    .A2(ld),
    .B(n_12860_o_0),
    .Y(n_12861_o_0));
 NAND2xp33_ASAP7_75t_R n_12862 (.A(ld),
    .B(text_in[124]),
    .Y(n_12862_o_0));
 OAI21xp33_ASAP7_75t_R n_12863 (.A1(_00652_),
    .A2(ld),
    .B(n_12862_o_0),
    .Y(n_12863_o_0));
 NAND2xp33_ASAP7_75t_R n_12864 (.A(ld),
    .B(text_in[125]),
    .Y(n_12864_o_0));
 OAI21xp33_ASAP7_75t_R n_12865 (.A1(_00651_),
    .A2(ld),
    .B(n_12864_o_0),
    .Y(n_12865_o_0));
 NAND2xp33_ASAP7_75t_R n_12866 (.A(ld),
    .B(text_in[126]),
    .Y(n_12866_o_0));
 OAI21xp33_ASAP7_75t_R n_12867 (.A1(_00650_),
    .A2(ld),
    .B(n_12866_o_0),
    .Y(n_12867_o_0));
 NAND2xp33_ASAP7_75t_R n_12868 (.A(ld),
    .B(text_in[127]),
    .Y(n_12868_o_0));
 OAI21xp33_ASAP7_75t_R n_12869 (.A1(_00649_),
    .A2(ld),
    .B(n_12868_o_0),
    .Y(n_12869_o_0));
 NAND2xp33_ASAP7_75t_R n_1287 (.A(n_889_o_0),
    .B(n_1121_o_0),
    .Y(n_1287_o_0));
 NAND2xp33_ASAP7_75t_R n_12870 (.A(_00647_),
    .B(_00648_),
    .Y(n_12870_o_0));
 OAI31xp33_ASAP7_75t_R n_12871 (.A1(n_12238_o_0),
    .A2(n_12870_o_0),
    .A3(n_12240_o_0),
    .B(rst),
    .Y(n_12871_o_0));
 INVx1_ASAP7_75t_R n_12872 (.A(_00648_),
    .Y(n_12872_o_0));
 INVx1_ASAP7_75t_R n_12873 (.A(rst),
    .Y(n_12873_o_0));
 OAI22xp33_ASAP7_75t_R n_12874 (.A1(n_12871_o_0),
    .A2(n_12872_o_0),
    .B1(n_827_o_0),
    .B2(n_12873_o_0),
    .Y(n_12874_o_0));
 AOI21xp33_ASAP7_75t_R n_12875 (.A1(_00645_),
    .A2(_00729_),
    .B(n_12870_o_0),
    .Y(n_12875_o_0));
 AOI21xp33_ASAP7_75t_R n_12876 (.A1(n_12239_o_0),
    .A2(n_12872_o_0),
    .B(n_12875_o_0),
    .Y(n_12876_o_0));
 AOI21xp33_ASAP7_75t_R n_12877 (.A1(n_827_o_0),
    .A2(n_12876_o_0),
    .B(n_12873_o_0),
    .Y(n_12877_o_0));
 OAI211xp5_ASAP7_75t_R n_12878 (.A1(n_12870_o_0),
    .A2(n_12238_o_0),
    .B(n_12240_o_0),
    .C(rst),
    .Y(n_12878_o_0));
 OAI21xp33_ASAP7_75t_R n_12879 (.A1(n_827_o_0),
    .A2(n_12873_o_0),
    .B(n_12878_o_0),
    .Y(n_12879_o_0));
 NAND2xp33_ASAP7_75t_R n_1288 (.A(n_864_o_0),
    .B(n_836_o_0),
    .Y(n_1288_o_0));
 XNOR2xp5_ASAP7_75t_R n_12880 (.A(_00645_),
    .B(n_12870_o_0),
    .Y(n_12880_o_0));
 NOR3xp33_ASAP7_75t_R n_12881 (.A(n_12880_o_0),
    .B(n_12871_o_0),
    .C(ld),
    .Y(n_12881_o_0));
 INVx1_ASAP7_75t_R n_12882 (.A(\u0/r0/rcnt_next[0] ),
    .Y(n_12882_o_0));
 NOR2xp33_ASAP7_75t_R n_12883 (.A(ld),
    .B(n_12882_o_0),
    .Y(n_12883_o_0));
 XNOR2xp5_ASAP7_75t_R n_12884 (.A(_11695_),
    .B(\u0/r0/rcnt_next[0] ),
    .Y(n_12884_o_0));
 NOR2xp33_ASAP7_75t_R n_12885 (.A(ld),
    .B(n_12884_o_0),
    .Y(n_12885_o_0));
 NOR2xp33_ASAP7_75t_R n_12886 (.A(_11695_),
    .B(\u0/r0/rcnt_next[0] ),
    .Y(n_12886_o_0));
 XOR2xp5_ASAP7_75t_R n_12887 (.A(_00644_),
    .B(n_12886_o_0),
    .Y(n_12887_o_0));
 NOR2xp33_ASAP7_75t_R n_12888 (.A(ld),
    .B(n_12887_o_0),
    .Y(n_12888_o_0));
 NOR3xp33_ASAP7_75t_R n_12889 (.A(_00644_),
    .B(_11695_),
    .C(\u0/r0/rcnt_next[0] ),
    .Y(n_12889_o_0));
 OAI21xp33_ASAP7_75t_R n_1289 (.A1(n_864_o_0),
    .A2(net32),
    .B(n_1288_o_0),
    .Y(n_1289_o_0));
 XOR2xp5_ASAP7_75t_R n_12890 (.A(_00859_),
    .B(n_12889_o_0),
    .Y(n_12890_o_0));
 NOR2xp33_ASAP7_75t_R n_12891 (.A(ld),
    .B(n_12890_o_0),
    .Y(n_12891_o_0));
 XNOR2xp5_ASAP7_75t_R n_12892 (.A(_00644_),
    .B(n_12886_o_0),
    .Y(n_12892_o_0));
 OAI31xp33_ASAP7_75t_R n_12893 (.A1(_11695_),
    .A2(n_12892_o_0),
    .A3(\u0/r0/rcnt_next[0] ),
    .B(n_827_o_0),
    .Y(n_12893_o_0));
 NOR2xp33_ASAP7_75t_R n_12894 (.A(n_12892_o_0),
    .B(n_12890_o_0),
    .Y(n_12894_o_0));
 NAND2xp33_ASAP7_75t_R n_12895 (.A(n_12884_o_0),
    .B(n_12894_o_0),
    .Y(n_12895_o_0));
 AND2x2_ASAP7_75t_R n_12896 (.A(n_12887_o_0),
    .B(n_12890_o_0),
    .Y(n_12896_o_0));
 NAND3xp33_ASAP7_75t_R n_12897 (.A(n_12896_o_0),
    .B(\u0/r0/rcnt_next[0] ),
    .C(_11695_),
    .Y(n_12897_o_0));
 AOI21xp33_ASAP7_75t_R n_12898 (.A1(n_12895_o_0),
    .A2(n_12897_o_0),
    .B(ld),
    .Y(n_12898_o_0));
 INVx1_ASAP7_75t_R n_12899 (.A(n_12894_o_0),
    .Y(n_12899_o_0));
 AOI211xp5_ASAP7_75t_R n_1290 (.A1(n_1289_o_0),
    .A2(n_878_o_0),
    .B(n_1209_o_0),
    .C(n_829_o_0),
    .Y(n_1290_o_0));
 OAI21xp33_ASAP7_75t_R n_12900 (.A1(\u0/r0/rcnt_next[0] ),
    .A2(n_12896_o_0),
    .B(_11695_),
    .Y(n_12900_o_0));
 AOI311xp33_ASAP7_75t_R n_12901 (.A1(n_12899_o_0),
    .A2(\u0/r0/rcnt_next[0] ),
    .A3(_11695_),
    .B(ld),
    .C(n_12900_o_0),
    .Y(n_12901_o_0));
 NAND2xp33_ASAP7_75t_R n_12902 (.A(n_12887_o_0),
    .B(n_12890_o_0),
    .Y(n_12902_o_0));
 NAND3xp33_ASAP7_75t_R n_12903 (.A(n_12902_o_0),
    .B(n_12887_o_0),
    .C(n_12886_o_0),
    .Y(n_12903_o_0));
 INVx1_ASAP7_75t_R n_12904 (.A(_11695_),
    .Y(n_12904_o_0));
 NAND3xp33_ASAP7_75t_R n_12905 (.A(n_12896_o_0),
    .B(n_12904_o_0),
    .C(\u0/r0/rcnt_next[0] ),
    .Y(n_12905_o_0));
 AOI21xp33_ASAP7_75t_R n_12906 (.A1(n_12903_o_0),
    .A2(n_12905_o_0),
    .B(ld),
    .Y(n_12906_o_0));
 AND3x1_ASAP7_75t_R n_12907 (.A(n_12894_o_0),
    .B(n_12884_o_0),
    .C(n_827_o_0),
    .Y(n_12907_o_0));
 AOI31xp33_ASAP7_75t_R n_12908 (.A1(n_12886_o_0),
    .A2(n_12888_o_0),
    .A3(n_12890_o_0),
    .B(n_12907_o_0),
    .Y(n_12908_o_0));
 INVx1_ASAP7_75t_R n_12909 (.A(n_12908_o_0),
    .Y(n_12909_o_0));
 AOI21xp33_ASAP7_75t_R n_1291 (.A1(n_1043_o_0),
    .A2(n_1287_o_0),
    .B(n_1290_o_0),
    .Y(n_1291_o_0));
 OAI21xp33_ASAP7_75t_R n_12910 (.A1(n_12887_o_0),
    .A2(n_12890_o_0),
    .B(n_12902_o_0),
    .Y(n_12910_o_0));
 NOR4xp25_ASAP7_75t_R n_12911 (.A(n_12910_o_0),
    .B(n_12882_o_0),
    .C(n_12904_o_0),
    .D(ld),
    .Y(n_12911_o_0));
 NAND3xp33_ASAP7_75t_R n_12912 (.A(n_12890_o_0),
    .B(n_827_o_0),
    .C(n_12892_o_0),
    .Y(n_12912_o_0));
 NOR3xp33_ASAP7_75t_R n_12913 (.A(n_12912_o_0),
    .B(n_12904_o_0),
    .C(\u0/r0/rcnt_next[0] ),
    .Y(n_12913_o_0));
 NOR3xp33_ASAP7_75t_R n_12914 (.A(n_12912_o_0),
    .B(n_12882_o_0),
    .C(_11695_),
    .Y(n_12914_o_0));
 XOR2xp5_ASAP7_75t_R n_12915 (.A(_11695_),
    .B(\u0/r0/rcnt_next[0] ),
    .Y(n_12915_o_0));
 INVx1_ASAP7_75t_R n_12916 (.A(n_909_o_1),
    .Y(n_12916_o_0));
 AO21x1_ASAP7_75t_R n_12917 (.A1(n_859_o_0),
    .A2(net32),
    .B(n_1229_o_0),
    .Y(n_12917_o_0));
 NAND2xp33_ASAP7_75t_R n_12918 (.A(n_1387_o_0),
    .B(n_1404_o_0),
    .Y(n_12918_o_0));
 OAI21xp33_ASAP7_75t_R n_12919 (.A1(n_1387_o_0),
    .A2(n_1404_o_0),
    .B(n_12918_o_0),
    .Y(n_12919_o_0));
 OAI22xp33_ASAP7_75t_R n_1292 (.A1(n_1285_o_0),
    .A2(n_1286_o_0),
    .B1(n_903_o_0),
    .B2(n_1291_o_0),
    .Y(n_1292_o_0));
 NAND2xp33_ASAP7_75t_R n_12920 (.A(n_1555_o_0),
    .B(n_1788_o_0),
    .Y(n_12920_o_0));
 NAND2xp33_ASAP7_75t_R n_12921 (.A(net99),
    .B(n_1380_o_0),
    .Y(n_12921_o_0));
 OAI21xp33_ASAP7_75t_R n_12922 (.A1(n_1380_o_0),
    .A2(net99),
    .B(n_12921_o_0),
    .Y(n_12922_o_0));
 NAND2xp33_ASAP7_75t_R n_12923 (.A(n_1912_o_0),
    .B(n_1916_o_0),
    .Y(n_12923_o_0));
 OAI21xp33_ASAP7_75t_R n_12924 (.A1(n_1916_o_0),
    .A2(n_1912_o_0),
    .B(n_12923_o_0),
    .Y(n_12924_o_0));
 NAND2xp33_ASAP7_75t_R n_12925 (.A(n_2075_o_0),
    .B(n_2314_o_0),
    .Y(n_12925_o_0));
 NAND2xp33_ASAP7_75t_R n_12926 (.A(n_1941_o_0),
    .B(n_1898_o_0),
    .Y(n_12926_o_0));
 OAI21xp33_ASAP7_75t_R n_12927 (.A1(n_1941_o_0),
    .A2(n_1898_o_0),
    .B(n_12926_o_0),
    .Y(n_12927_o_0));
 XNOR2xp5_ASAP7_75t_R n_12928 (.A(n_2505_o_0),
    .B(net102),
    .Y(n_12928_o_0));
 INVx1_ASAP7_75t_R n_12929 (.A(n_2920_o_0),
    .Y(n_12929_o_0));
 AOI21xp33_ASAP7_75t_R n_1293 (.A1(n_971_o_0),
    .A2(n_1292_o_0),
    .B(n_931_o_0),
    .Y(n_1293_o_0));
 OAI21xp33_ASAP7_75t_R n_12930 (.A1(n_2505_o_0),
    .A2(net101),
    .B(n_2836_o_0),
    .Y(n_12930_o_0));
 OAI21xp33_ASAP7_75t_R n_12931 (.A1(n_3125_o_0),
    .A2(n_3124_o_0),
    .B(n_3540_o_0),
    .Y(n_12931_o_0));
 NAND2xp33_ASAP7_75t_R n_12932 (.A(net40),
    .B(net36),
    .Y(n_12932_o_0));
 OAI21xp33_ASAP7_75t_R n_12933 (.A1(net40),
    .A2(net36),
    .B(n_12932_o_0),
    .Y(n_12933_o_0));
 OAI33xp33_ASAP7_75t_R n_12934 (.A1(n_3734_o_0),
    .A2(net30),
    .A3(n_3672_o_0),
    .B1(n_3658_o_0),
    .B2(n_3707_o_0),
    .B3(net25),
    .Y(n_12934_o_0));
 OAI33xp33_ASAP7_75t_R n_12935 (.A1(n_3658_o_0),
    .A2(n_3707_o_0),
    .A3(net72),
    .B1(net30),
    .B2(n_3709_o_0),
    .B3(n_3682_o_0),
    .Y(n_12935_o_0));
 XNOR2xp5_ASAP7_75t_R n_12936 (.A(net82),
    .B(n_4287_o_0),
    .Y(n_12936_o_0));
 OAI21xp33_ASAP7_75t_R n_12937 (.A1(net47),
    .A2(net59),
    .B(n_4327_o_0),
    .Y(n_12937_o_0));
 NAND2xp33_ASAP7_75t_R n_12938 (.A(n_4752_o_0),
    .B(n_4751_o_0),
    .Y(n_12938_o_0));
 OAI33xp33_ASAP7_75t_R n_12939 (.A1(n_4999_o_0),
    .A2(n_4974_o_0),
    .A3(n_4899_o_0),
    .B1(n_4949_o_0),
    .B2(net69),
    .B3(n_4898_o_0),
    .Y(n_12939_o_0));
 OAI21xp33_ASAP7_75t_R n_1294 (.A1(n_971_o_0),
    .A2(n_1283_o_0),
    .B(n_1293_o_0),
    .Y(n_1294_o_0));
 OAI33xp33_ASAP7_75t_R n_12940 (.A1(net60),
    .A2(n_4999_o_0),
    .A3(n_4974_o_0),
    .B1(n_5019_o_0),
    .B2(net69),
    .B3(n_4872_o_0),
    .Y(n_12940_o_0));
 INVx1_ASAP7_75t_R n_12941 (.A(n_5378_o_0),
    .Y(n_12941_o_0));
 NAND2xp33_ASAP7_75t_R n_12942 (.A(n_5484_o_0),
    .B(n_5459_o_0),
    .Y(n_12942_o_0));
 OAI21xp33_ASAP7_75t_R n_12943 (.A1(n_5484_o_0),
    .A2(n_5459_o_0),
    .B(n_12942_o_0),
    .Y(n_12943_o_0));
 OAI33xp33_ASAP7_75t_R n_12944 (.A1(n_5529_o_0),
    .A2(n_5573_o_0),
    .A3(net54),
    .B1(n_5469_o_0),
    .B2(n_5549_o_0),
    .B3(n_5467_o_0),
    .Y(n_12944_o_0));
 OAI21xp33_ASAP7_75t_R n_12945 (.A1(n_6030_o_0),
    .A2(n_6017_o_0),
    .B(n_6052_o_0),
    .Y(n_12945_o_0));
 OAI21xp33_ASAP7_75t_R n_12946 (.A1(n_6039_o_0),
    .A2(n_6062_o_0),
    .B(n_6278_o_0),
    .Y(n_12946_o_0));
 NAND2xp33_ASAP7_75t_R n_12947 (.A(n_6405_o_0),
    .B(n_6215_o_0),
    .Y(n_12947_o_0));
 OAI21xp33_ASAP7_75t_R n_12948 (.A1(n_6601_o_0),
    .A2(n_6588_o_0),
    .B(n_6862_o_0),
    .Y(n_12948_o_0));
 INVx1_ASAP7_75t_R n_12949 (.A(n_7062_o_0),
    .Y(n_12949_o_0));
 OAI31xp33_ASAP7_75t_R n_1295 (.A1(n_1264_o_0),
    .A2(n_1274_o_0),
    .A3(n_930_o_0),
    .B(n_1294_o_0),
    .Y(n_1295_o_0));
 OAI21xp33_ASAP7_75t_R n_12950 (.A1(net79),
    .A2(n_7182_o_0),
    .B(n_7303_o_0),
    .Y(n_12950_o_0));
 AO21x1_ASAP7_75t_R n_12951 (.A1(n_7201_o_0),
    .A2(net46),
    .B(n_7263_o_0),
    .Y(n_12951_o_0));
 NAND2xp33_ASAP7_75t_R n_12952 (.A(net34),
    .B(n_7768_o_0),
    .Y(n_12952_o_0));
 OAI21xp33_ASAP7_75t_R n_12953 (.A1(n_7768_o_0),
    .A2(net34),
    .B(n_12952_o_0),
    .Y(n_12953_o_0));
 OAI21xp33_ASAP7_75t_R n_12954 (.A1(n_7796_o_0),
    .A2(net34),
    .B(n_7944_o_0),
    .Y(n_12954_o_0));
 NAND2xp33_ASAP7_75t_R n_12955 (.A(net67),
    .B(net38),
    .Y(n_12955_o_0));
 OAI21xp33_ASAP7_75t_R n_12956 (.A1(net67),
    .A2(net38),
    .B(n_12955_o_0),
    .Y(n_12956_o_0));
 OAI21xp33_ASAP7_75t_R n_12957 (.A1(net73),
    .A2(net38),
    .B(n_8679_o_0),
    .Y(n_12957_o_0));
 NAND2xp33_ASAP7_75t_R n_12958 (.A(net19),
    .B(n_8915_o_0),
    .Y(n_12958_o_0));
 OAI21xp33_ASAP7_75t_R n_12959 (.A1(n_8915_o_0),
    .A2(net19),
    .B(n_12958_o_0),
    .Y(n_12959_o_0));
 NOR3xp33_ASAP7_75t_R n_1296 (.A(n_878_o_0),
    .B(n_913_o_0),
    .C(n_881_o_0),
    .Y(n_1296_o_0));
 AO21x1_ASAP7_75t_R n_12960 (.A1(net19),
    .A2(n_8947_o_0),
    .B(n_9197_o_0),
    .Y(n_12960_o_0));
 NAND2xp33_ASAP7_75t_R n_12961 (.A(n_9451_o_0),
    .B(net26),
    .Y(n_12961_o_0));
 OAI21xp33_ASAP7_75t_R n_12962 (.A1(n_9451_o_0),
    .A2(net26),
    .B(n_12961_o_0),
    .Y(n_12962_o_0));
 NAND2xp33_ASAP7_75t_R n_12963 (.A(net26),
    .B(n_9435_o_0),
    .Y(n_12963_o_0));
 OAI21xp33_ASAP7_75t_R n_12964 (.A1(n_9435_o_0),
    .A2(net26),
    .B(n_12963_o_0),
    .Y(n_12964_o_0));
 OAI33xp33_ASAP7_75t_R n_12965 (.A1(net24),
    .A2(n_10019_o_0),
    .A3(n_10023_o_0),
    .B1(n_10074_o_0),
    .B2(n_10024_o_0),
    .B3(n_10011_o_0),
    .Y(n_12965_o_0));
 NAND2xp33_ASAP7_75t_R n_12966 (.A(net56),
    .B(n_10043_o_0),
    .Y(n_12966_o_0));
 OAI21xp33_ASAP7_75t_R n_12967 (.A1(net56),
    .A2(n_10043_o_0),
    .B(n_12966_o_0),
    .Y(n_12967_o_0));
 INVx1_ASAP7_75t_R n_12968 (.A(n_10488_o_0),
    .Y(n_12968_o_0));
 OAI33xp33_ASAP7_75t_R n_12969 (.A1(n_10591_o_0),
    .A2(n_10562_o_0),
    .A3(n_10566_o_0),
    .B1(n_10652_o_0),
    .B2(n_10567_o_0),
    .B3(n_10590_o_0),
    .Y(n_12969_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_1297 (.A1(n_881_o_0),
    .A2(n_889_o_0),
    .B(n_866_o_0),
    .C(n_878_o_0),
    .D(n_1296_o_0),
    .Y(n_1297_o_0));
 OAI33xp33_ASAP7_75t_R n_12970 (.A1(net43),
    .A2(n_10562_o_0),
    .A3(n_10566_o_0),
    .B1(n_10579_o_0),
    .B2(n_10567_o_0),
    .B3(n_10668_o_0),
    .Y(n_12970_o_0));
 NAND2xp33_ASAP7_75t_R n_12971 (.A(net58),
    .B(net35),
    .Y(n_12971_o_0));
 OAI21xp33_ASAP7_75t_R n_12972 (.A1(net58),
    .A2(net35),
    .B(n_12971_o_0),
    .Y(n_12972_o_0));
 NAND2xp33_ASAP7_75t_R n_12973 (.A(n_11503_o_0),
    .B(n_11532_o_0),
    .Y(n_12973_o_0));
 OAI21xp33_ASAP7_75t_R n_12974 (.A1(n_11733_o_0),
    .A2(n_11707_o_0),
    .B(n_11923_o_0),
    .Y(n_12974_o_0));
 INVx1_ASAP7_75t_R n_12975 (.A(_00646_),
    .Y(n_12975_o_0));
 INVx1_ASAP7_75t_R n_12976 (.A(_00730_),
    .Y(n_12976_o_0));
 INVx1_ASAP7_75t_R n_12977 (.A(_00758_),
    .Y(n_12977_o_0));
 INVx1_ASAP7_75t_R n_12978 (.A(_00759_),
    .Y(n_12978_o_0));
 INVx1_ASAP7_75t_R n_12979 (.A(_00760_),
    .Y(n_12979_o_0));
 AOI211xp5_ASAP7_75t_R n_1298 (.A1(n_1028_o_0),
    .A2(n_957_o_0),
    .B(n_1152_o_0),
    .C(n_891_o_0),
    .Y(n_1298_o_0));
 INVx1_ASAP7_75t_R n_12980 (.A(_00761_),
    .Y(n_12980_o_0));
 INVx1_ASAP7_75t_R n_12981 (.A(_00786_),
    .Y(n_12981_o_0));
 INVx1_ASAP7_75t_R n_12982 (.A(_00787_),
    .Y(n_12982_o_0));
 INVx1_ASAP7_75t_R n_12983 (.A(_00788_),
    .Y(n_12983_o_0));
 INVx1_ASAP7_75t_R n_12984 (.A(_00789_),
    .Y(n_12984_o_0));
 INVx1_ASAP7_75t_R n_12985 (.A(_00790_),
    .Y(n_12985_o_0));
 INVx1_ASAP7_75t_R n_12986 (.A(_00791_),
    .Y(n_12986_o_0));
 INVx1_ASAP7_75t_R n_12987 (.A(_00764_),
    .Y(n_12987_o_0));
 INVx1_ASAP7_75t_R n_12988 (.A(_00792_),
    .Y(n_12988_o_0));
 INVx1_ASAP7_75t_R n_12989 (.A(_00793_),
    .Y(n_12989_o_0));
 AOI31xp33_ASAP7_75t_R n_1299 (.A1(n_891_o_0),
    .A2(n_1189_o_0),
    .A3(n_1297_o_0),
    .B(n_1298_o_0),
    .Y(n_1299_o_0));
 INVx1_ASAP7_75t_R n_12990 (.A(_00818_),
    .Y(n_12990_o_0));
 INVx1_ASAP7_75t_R n_12991 (.A(_00819_),
    .Y(n_12991_o_0));
 INVx1_ASAP7_75t_R n_12992 (.A(_00820_),
    .Y(n_12992_o_0));
 INVx1_ASAP7_75t_R n_12993 (.A(_00821_),
    .Y(n_12993_o_0));
 INVx1_ASAP7_75t_R n_12994 (.A(_00822_),
    .Y(n_12994_o_0));
 INVx1_ASAP7_75t_R n_12995 (.A(_00823_),
    .Y(n_12995_o_0));
 INVx1_ASAP7_75t_R n_12996 (.A(_00824_),
    .Y(n_12996_o_0));
 INVx1_ASAP7_75t_R n_12997 (.A(_00825_),
    .Y(n_12997_o_0));
 INVx1_ASAP7_75t_R n_12998 (.A(_00765_),
    .Y(n_12998_o_0));
 INVx1_ASAP7_75t_R n_12999 (.A(_00850_),
    .Y(n_12999_o_0));
 AOI211xp5_ASAP7_75t_R n_1300 (.A1(n_877_o_0),
    .A2(n_933_o_0),
    .B(n_881_o_0),
    .C(n_864_o_0),
    .Y(n_1300_o_0));
 INVx1_ASAP7_75t_R n_13000 (.A(_00851_),
    .Y(n_13000_o_0));
 INVx1_ASAP7_75t_R n_13001 (.A(_00852_),
    .Y(n_13001_o_0));
 INVx1_ASAP7_75t_R n_13002 (.A(_00853_),
    .Y(n_13002_o_0));
 INVx1_ASAP7_75t_R n_13003 (.A(_00854_),
    .Y(n_13003_o_0));
 INVx1_ASAP7_75t_R n_13004 (.A(_00855_),
    .Y(n_13004_o_0));
 INVx1_ASAP7_75t_R n_13005 (.A(_00856_),
    .Y(n_13005_o_0));
 INVx1_ASAP7_75t_R n_13006 (.A(_00857_),
    .Y(n_13006_o_0));
 INVx1_ASAP7_75t_R n_13007 (.A(_00766_),
    .Y(n_13007_o_0));
 INVx1_ASAP7_75t_R n_13008 (.A(_00767_),
    .Y(n_13008_o_0));
 INVx1_ASAP7_75t_R n_13009 (.A(_00768_),
    .Y(n_13009_o_0));
 NOR3xp33_ASAP7_75t_R n_1301 (.A(n_996_o_0),
    .B(n_1300_o_0),
    .C(n_829_o_0),
    .Y(n_1301_o_0));
 INVx1_ASAP7_75t_R n_13010 (.A(_00769_),
    .Y(n_13010_o_0));
 INVx1_ASAP7_75t_R n_13011 (.A(_00794_),
    .Y(n_13011_o_0));
 INVx1_ASAP7_75t_R n_13012 (.A(_00795_),
    .Y(n_13012_o_0));
 INVx1_ASAP7_75t_R n_13013 (.A(_00796_),
    .Y(n_13013_o_0));
 INVx1_ASAP7_75t_R n_13014 (.A(_00797_),
    .Y(n_13014_o_0));
 INVx1_ASAP7_75t_R n_13015 (.A(_00731_),
    .Y(n_13015_o_0));
 INVx1_ASAP7_75t_R n_13016 (.A(_00798_),
    .Y(n_13016_o_0));
 INVx1_ASAP7_75t_R n_13017 (.A(_00799_),
    .Y(n_13017_o_0));
 INVx1_ASAP7_75t_R n_13018 (.A(_00800_),
    .Y(n_13018_o_0));
 INVx1_ASAP7_75t_R n_13019 (.A(_00801_),
    .Y(n_13019_o_0));
 OAI21xp33_ASAP7_75t_R n_1302 (.A1(n_935_o_0),
    .A2(n_878_o_0),
    .B(n_829_o_0),
    .Y(n_1302_o_0));
 INVx1_ASAP7_75t_R n_13020 (.A(_00826_),
    .Y(n_13020_o_0));
 INVx1_ASAP7_75t_R n_13021 (.A(_00827_),
    .Y(n_13021_o_0));
 INVx1_ASAP7_75t_R n_13022 (.A(_00828_),
    .Y(n_13022_o_0));
 INVx1_ASAP7_75t_R n_13023 (.A(_00829_),
    .Y(n_13023_o_0));
 INVx1_ASAP7_75t_R n_13024 (.A(_00830_),
    .Y(n_13024_o_0));
 INVx1_ASAP7_75t_R n_13025 (.A(_00831_),
    .Y(n_13025_o_0));
 INVx1_ASAP7_75t_R n_13026 (.A(_00732_),
    .Y(n_13026_o_0));
 INVx1_ASAP7_75t_R n_13027 (.A(_00832_),
    .Y(n_13027_o_0));
 INVx1_ASAP7_75t_R n_13028 (.A(_00833_),
    .Y(n_13028_o_0));
 INVx1_ASAP7_75t_R n_13029 (.A(_00738_),
    .Y(n_13029_o_0));
 AOI21xp33_ASAP7_75t_R n_1303 (.A1(n_878_o_0),
    .A2(n_1181_o_0),
    .B(n_1302_o_0),
    .Y(n_1303_o_0));
 INVx1_ASAP7_75t_R n_13030 (.A(_00739_),
    .Y(n_13030_o_0));
 INVx1_ASAP7_75t_R n_13031 (.A(_00740_),
    .Y(n_13031_o_0));
 INVx1_ASAP7_75t_R n_13032 (.A(_00741_),
    .Y(n_13032_o_0));
 INVx1_ASAP7_75t_R n_13033 (.A(_00742_),
    .Y(n_13033_o_0));
 INVx1_ASAP7_75t_R n_13034 (.A(_00743_),
    .Y(n_13034_o_0));
 INVx1_ASAP7_75t_R n_13035 (.A(_00744_),
    .Y(n_13035_o_0));
 INVx1_ASAP7_75t_R n_13036 (.A(_00745_),
    .Y(n_13036_o_0));
 INVx1_ASAP7_75t_R n_13037 (.A(_00733_),
    .Y(n_13037_o_0));
 INVx1_ASAP7_75t_R n_13038 (.A(_00770_),
    .Y(n_13038_o_0));
 INVx1_ASAP7_75t_R n_13039 (.A(_00771_),
    .Y(n_13039_o_0));
 NOR3xp33_ASAP7_75t_R n_1304 (.A(n_1301_o_0),
    .B(n_1303_o_0),
    .C(n_904_o_0),
    .Y(n_1304_o_0));
 INVx1_ASAP7_75t_R n_13040 (.A(_00772_),
    .Y(n_13040_o_0));
 INVx1_ASAP7_75t_R n_13041 (.A(_00773_),
    .Y(n_13041_o_0));
 INVx1_ASAP7_75t_R n_13042 (.A(_00774_),
    .Y(n_13042_o_0));
 INVx1_ASAP7_75t_R n_13043 (.A(_00775_),
    .Y(n_13043_o_0));
 INVx1_ASAP7_75t_R n_13044 (.A(_00776_),
    .Y(n_13044_o_0));
 INVx1_ASAP7_75t_R n_13045 (.A(_00777_),
    .Y(n_13045_o_0));
 INVx1_ASAP7_75t_R n_13046 (.A(_00802_),
    .Y(n_13046_o_0));
 INVx1_ASAP7_75t_R n_13047 (.A(_00803_),
    .Y(n_13047_o_0));
 INVx1_ASAP7_75t_R n_13048 (.A(_00734_),
    .Y(n_13048_o_0));
 INVx1_ASAP7_75t_R n_13049 (.A(_00804_),
    .Y(n_13049_o_0));
 AOI21xp33_ASAP7_75t_R n_1305 (.A1(n_904_o_0),
    .A2(n_1299_o_0),
    .B(n_1304_o_0),
    .Y(n_1305_o_0));
 INVx1_ASAP7_75t_R n_13050 (.A(_00805_),
    .Y(n_13050_o_0));
 INVx1_ASAP7_75t_R n_13051 (.A(_00806_),
    .Y(n_13051_o_0));
 INVx1_ASAP7_75t_R n_13052 (.A(_00807_),
    .Y(n_13052_o_0));
 INVx1_ASAP7_75t_R n_13053 (.A(_00808_),
    .Y(n_13053_o_0));
 INVx1_ASAP7_75t_R n_13054 (.A(_00809_),
    .Y(n_13054_o_0));
 INVx1_ASAP7_75t_R n_13055 (.A(_00834_),
    .Y(n_13055_o_0));
 INVx1_ASAP7_75t_R n_13056 (.A(_00835_),
    .Y(n_13056_o_0));
 INVx1_ASAP7_75t_R n_13057 (.A(_00836_),
    .Y(n_13057_o_0));
 INVx1_ASAP7_75t_R n_13058 (.A(_00837_),
    .Y(n_13058_o_0));
 INVx1_ASAP7_75t_R n_13059 (.A(_00735_),
    .Y(n_13059_o_0));
 NAND3xp33_ASAP7_75t_R n_1306 (.A(n_882_o_0),
    .B(n_990_o_0),
    .C(n_878_o_0),
    .Y(n_1306_o_0));
 INVx1_ASAP7_75t_R n_13060 (.A(_00838_),
    .Y(n_13060_o_0));
 INVx1_ASAP7_75t_R n_13061 (.A(_00839_),
    .Y(n_13061_o_0));
 INVx1_ASAP7_75t_R n_13062 (.A(_00840_),
    .Y(n_13062_o_0));
 INVx1_ASAP7_75t_R n_13063 (.A(_00841_),
    .Y(n_13063_o_0));
 INVx1_ASAP7_75t_R n_13064 (.A(_00746_),
    .Y(n_13064_o_0));
 INVx1_ASAP7_75t_R n_13065 (.A(_00747_),
    .Y(n_13065_o_0));
 INVx1_ASAP7_75t_R n_13066 (.A(_00748_),
    .Y(n_13066_o_0));
 INVx1_ASAP7_75t_R n_13067 (.A(_00749_),
    .Y(n_13067_o_0));
 INVx1_ASAP7_75t_R n_13068 (.A(_00750_),
    .Y(n_13068_o_0));
 INVx1_ASAP7_75t_R n_13069 (.A(_00751_),
    .Y(n_13069_o_0));
 OAI31xp33_ASAP7_75t_R n_1307 (.A1(n_878_o_0),
    .A2(n_989_o_0),
    .A3(n_994_o_0),
    .B(n_1306_o_0),
    .Y(n_1307_o_0));
 INVx1_ASAP7_75t_R n_13070 (.A(_00736_),
    .Y(n_13070_o_0));
 INVx1_ASAP7_75t_R n_13071 (.A(_00752_),
    .Y(n_13071_o_0));
 INVx1_ASAP7_75t_R n_13072 (.A(_00753_),
    .Y(n_13072_o_0));
 INVx1_ASAP7_75t_R n_13073 (.A(_00778_),
    .Y(n_13073_o_0));
 INVx1_ASAP7_75t_R n_13074 (.A(_00779_),
    .Y(n_13074_o_0));
 INVx1_ASAP7_75t_R n_13075 (.A(_00780_),
    .Y(n_13075_o_0));
 INVx1_ASAP7_75t_R n_13076 (.A(_00781_),
    .Y(n_13076_o_0));
 INVx1_ASAP7_75t_R n_13077 (.A(_00782_),
    .Y(n_13077_o_0));
 INVx1_ASAP7_75t_R n_13078 (.A(_00783_),
    .Y(n_13078_o_0));
 INVx1_ASAP7_75t_R n_13079 (.A(_00784_),
    .Y(n_13079_o_0));
 AOI211xp5_ASAP7_75t_R n_1308 (.A1(n_1246_o_0),
    .A2(n_886_o_0),
    .B(n_903_o_0),
    .C(n_1041_o_0),
    .Y(n_1308_o_0));
 INVx1_ASAP7_75t_R n_13080 (.A(_00785_),
    .Y(n_13080_o_0));
 INVx1_ASAP7_75t_R n_13081 (.A(_00737_),
    .Y(n_13081_o_0));
 INVx1_ASAP7_75t_R n_13082 (.A(_00810_),
    .Y(n_13082_o_0));
 INVx1_ASAP7_75t_R n_13083 (.A(_00811_),
    .Y(n_13083_o_0));
 INVx1_ASAP7_75t_R n_13084 (.A(_00812_),
    .Y(n_13084_o_0));
 INVx1_ASAP7_75t_R n_13085 (.A(_00813_),
    .Y(n_13085_o_0));
 INVx1_ASAP7_75t_R n_13086 (.A(_00814_),
    .Y(n_13086_o_0));
 INVx1_ASAP7_75t_R n_13087 (.A(_00815_),
    .Y(n_13087_o_0));
 INVx1_ASAP7_75t_R n_13088 (.A(_00816_),
    .Y(n_13088_o_0));
 INVx1_ASAP7_75t_R n_13089 (.A(_00817_),
    .Y(n_13089_o_0));
 AOI21xp33_ASAP7_75t_R n_1309 (.A1(n_903_o_0),
    .A2(n_1307_o_0),
    .B(n_1308_o_0),
    .Y(n_1309_o_0));
 INVx1_ASAP7_75t_R n_13090 (.A(_00842_),
    .Y(n_13090_o_0));
 INVx1_ASAP7_75t_R n_13091 (.A(_00843_),
    .Y(n_13091_o_0));
 INVx1_ASAP7_75t_R n_13092 (.A(_00762_),
    .Y(n_13092_o_0));
 INVx1_ASAP7_75t_R n_13093 (.A(_00844_),
    .Y(n_13093_o_0));
 INVx1_ASAP7_75t_R n_13094 (.A(_00845_),
    .Y(n_13094_o_0));
 INVx1_ASAP7_75t_R n_13095 (.A(_00846_),
    .Y(n_13095_o_0));
 INVx1_ASAP7_75t_R n_13096 (.A(_00847_),
    .Y(n_13096_o_0));
 INVx1_ASAP7_75t_R n_13097 (.A(_00848_),
    .Y(n_13097_o_0));
 INVx1_ASAP7_75t_R n_13098 (.A(_00849_),
    .Y(n_13098_o_0));
 INVx1_ASAP7_75t_R n_13099 (.A(_00754_),
    .Y(n_13099_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_1310 (.A1(n_847_o_0),
    .A2(n_859_o_0),
    .B(n_880_o_0),
    .C(net32),
    .D(n_878_o_0),
    .Y(n_1310_o_0));
 INVx1_ASAP7_75t_R n_13100 (.A(_00755_),
    .Y(n_13100_o_0));
 INVx1_ASAP7_75t_R n_13101 (.A(_00756_),
    .Y(n_13101_o_0));
 INVx1_ASAP7_75t_R n_13102 (.A(_00757_),
    .Y(n_13102_o_0));
 INVx1_ASAP7_75t_R n_13103 (.A(_00763_),
    .Y(n_13103_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1311 (.A1(n_878_o_0),
    .A2(n_956_o_0),
    .B(n_1310_o_0),
    .C(n_983_o_0),
    .Y(n_1311_o_0));
 AOI31xp33_ASAP7_75t_R n_1312 (.A1(n_836_o_0),
    .A2(n_860_o_0),
    .A3(n_877_o_0),
    .B(n_903_o_0),
    .Y(n_1312_o_0));
 OAI21xp33_ASAP7_75t_R n_1313 (.A1(n_877_o_0),
    .A2(n_913_o_0),
    .B(n_1312_o_0),
    .Y(n_1313_o_0));
 OAI21xp33_ASAP7_75t_R n_1314 (.A1(n_904_o_0),
    .A2(n_1311_o_0),
    .B(n_1313_o_0),
    .Y(n_1314_o_0));
 OAI21xp33_ASAP7_75t_R n_1315 (.A1(net42),
    .A2(n_1314_o_0),
    .B(n_930_o_0),
    .Y(n_1315_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1316 (.A1(n_1309_o_0),
    .A2(net42),
    .B(n_1315_o_0),
    .C(n_972_o_0),
    .Y(n_1316_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_1317 (.A1(key[22]),
    .A2(ld),
    .B(n_929_o_0),
    .C(n_1305_o_0),
    .D(n_1316_o_0),
    .Y(n_1317_o_0));
 INVx1_ASAP7_75t_R n_1318 (.A(n_1317_o_0),
    .Y(n_1318_o_0));
 AOI211xp5_ASAP7_75t_R n_1319 (.A1(n_889_o_0),
    .A2(n_881_o_0),
    .B(n_878_o_0),
    .C(n_1155_o_0),
    .Y(n_1319_o_0));
 OAI211xp5_ASAP7_75t_R n_1320 (.A1(n_1167_o_0),
    .A2(n_1006_o_0),
    .B(n_1102_o_0),
    .C(n_891_o_0),
    .Y(n_1320_o_0));
 OAI31xp33_ASAP7_75t_R n_1321 (.A1(n_1034_o_0),
    .A2(n_1319_o_0),
    .A3(net15),
    .B(n_1320_o_0),
    .Y(n_1321_o_0));
 AOI31xp33_ASAP7_75t_R n_1322 (.A1(n_891_o_0),
    .A2(n_1200_o_0),
    .A3(n_1167_o_0),
    .B(n_903_o_0),
    .Y(n_1322_o_0));
 AOI211xp5_ASAP7_75t_R n_1323 (.A1(n_861_o_0),
    .A2(n_878_o_0),
    .B(n_891_o_0),
    .C(n_1267_o_0),
    .Y(n_1323_o_0));
 OAI21xp33_ASAP7_75t_R n_1324 (.A1(n_995_o_0),
    .A2(n_945_o_0),
    .B(n_1323_o_0),
    .Y(n_1324_o_0));
 AOI21xp33_ASAP7_75t_R n_1325 (.A1(n_1322_o_0),
    .A2(n_1324_o_0),
    .B(n_930_o_0),
    .Y(n_1325_o_0));
 OAI21xp33_ASAP7_75t_R n_1326 (.A1(n_1321_o_0),
    .A2(n_904_o_0),
    .B(n_1325_o_0),
    .Y(n_1326_o_0));
 AOI21xp33_ASAP7_75t_R n_1327 (.A1(net32),
    .A2(n_913_o_0),
    .B(n_890_o_0),
    .Y(n_1327_o_0));
 OAI211xp5_ASAP7_75t_R n_1328 (.A1(n_1327_o_0),
    .A2(n_1166_o_0),
    .B(n_903_o_0),
    .C(net16),
    .Y(n_1328_o_0));
 OAI31xp33_ASAP7_75t_R n_1329 (.A1(n_907_o_0),
    .A2(n_1060_o_0),
    .A3(n_877_o_0),
    .B(n_1234_o_0),
    .Y(n_1329_o_0));
 OAI211xp5_ASAP7_75t_R n_1330 (.A1(n_957_o_0),
    .A2(n_881_o_0),
    .B(n_877_o_0),
    .C(n_953_o_0),
    .Y(n_1330_o_0));
 AOI31xp33_ASAP7_75t_R n_1331 (.A1(n_1330_o_0),
    .A2(n_1094_o_0),
    .A3(n_891_o_0),
    .B(n_903_o_0),
    .Y(n_1331_o_0));
 OAI21xp33_ASAP7_75t_R n_1332 (.A1(net14),
    .A2(n_1329_o_0),
    .B(n_1331_o_0),
    .Y(n_1332_o_0));
 NAND3xp33_ASAP7_75t_R n_1333 (.A(n_957_o_0),
    .B(n_881_o_0),
    .C(n_878_o_0),
    .Y(n_1333_o_0));
 OAI31xp33_ASAP7_75t_R n_1334 (.A1(n_878_o_0),
    .A2(net32),
    .A3(n_1044_o_0),
    .B(n_1333_o_0),
    .Y(n_1334_o_0));
 NAND3xp33_ASAP7_75t_R n_1335 (.A(n_1334_o_0),
    .B(n_903_o_0),
    .C(net14),
    .Y(n_1335_o_0));
 NAND4xp25_ASAP7_75t_R n_1336 (.A(n_1328_o_0),
    .B(n_1332_o_0),
    .C(n_1335_o_0),
    .D(n_930_o_0),
    .Y(n_1336_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1337 (.A1(n_1326_o_0),
    .A2(n_1336_o_0),
    .B(n_1317_o_0),
    .C(n_971_o_0),
    .Y(n_1337_o_0));
 OAI21xp33_ASAP7_75t_R n_1338 (.A1(n_1318_o_0),
    .A2(n_971_o_0),
    .B(n_1337_o_0),
    .Y(n_1338_o_0));
 XNOR2xp5_ASAP7_75t_R n_1339 (.A(_00438_),
    .B(_00875_),
    .Y(n_1339_o_0));
 INVx1_ASAP7_75t_R n_1340 (.A(n_1339_o_0),
    .Y(n_1340_o_0));
 XNOR2xp5_ASAP7_75t_R n_1341 (.A(_00907_),
    .B(n_1340_o_0),
    .Y(n_1341_o_0));
 INVx1_ASAP7_75t_R n_1342 (.A(_00939_),
    .Y(n_1342_o_0));
 NAND2xp33_ASAP7_75t_R n_1343 (.A(n_1342_o_0),
    .B(n_1341_o_0),
    .Y(n_1343_o_0));
 OAI21xp33_ASAP7_75t_R n_1344 (.A1(n_1341_o_0),
    .A2(n_1342_o_0),
    .B(n_1343_o_0),
    .Y(n_1344_o_0));
 XOR2xp5_ASAP7_75t_R n_1345 (.A(_00971_),
    .B(n_1344_o_0),
    .Y(n_1345_o_0));
 OR2x2_ASAP7_75t_R n_1346 (.A(key[15]),
    .B(n_827_o_0),
    .Y(n_1346_o_0));
 OAI21xp33_ASAP7_75t_R n_1347 (.A1(ld),
    .A2(n_1345_o_0),
    .B(n_1346_o_0),
    .Y(n_1347_o_0));
 XNOR2xp5_ASAP7_75t_R n_1348 (.A(_00437_),
    .B(_00874_),
    .Y(n_1348_o_0));
 NAND2xp33_ASAP7_75t_R n_1349 (.A(_00906_),
    .B(n_1348_o_0),
    .Y(n_1349_o_0));
 OAI21xp33_ASAP7_75t_R n_1350 (.A1(_00906_),
    .A2(n_1348_o_0),
    .B(n_1349_o_0),
    .Y(n_1350_o_0));
 NAND2xp33_ASAP7_75t_R n_1351 (.A(_00938_),
    .B(n_1350_o_0),
    .Y(n_1351_o_0));
 OAI21xp33_ASAP7_75t_R n_1352 (.A1(_00938_),
    .A2(n_1350_o_0),
    .B(n_1351_o_0),
    .Y(n_1352_o_0));
 NOR2xp33_ASAP7_75t_R n_1353 (.A(_00970_),
    .B(n_1352_o_0),
    .Y(n_1353_o_0));
 AOI211xp5_ASAP7_75t_R n_1354 (.A1(n_1352_o_0),
    .A2(_00970_),
    .B(n_1353_o_0),
    .C(ld),
    .Y(n_1354_o_0));
 AOI21xp33_ASAP7_75t_R n_1355 (.A1(key[14]),
    .A2(ld),
    .B(n_1354_o_0),
    .Y(n_1355_o_0));
 XOR2xp5_ASAP7_75t_R n_1356 (.A(_00435_),
    .B(_00872_),
    .Y(n_1356_o_0));
 XNOR2xp5_ASAP7_75t_R n_1357 (.A(_00904_),
    .B(n_1356_o_0),
    .Y(n_1357_o_0));
 XNOR2xp5_ASAP7_75t_R n_1358 (.A(_00936_),
    .B(n_1357_o_0),
    .Y(n_1358_o_0));
 INVx1_ASAP7_75t_R n_1359 (.A(_00968_),
    .Y(n_1359_o_0));
 NAND2xp33_ASAP7_75t_R n_1360 (.A(n_1359_o_0),
    .B(n_1358_o_0),
    .Y(n_1360_o_0));
 OAI21xp33_ASAP7_75t_R n_1361 (.A1(n_1358_o_0),
    .A2(n_1359_o_0),
    .B(n_1360_o_0),
    .Y(n_1361_o_0));
 NOR2xp33_ASAP7_75t_R n_1362 (.A(key[12]),
    .B(n_827_o_0),
    .Y(n_1362_o_0));
 AOI21x1_ASAP7_75t_R n_1363 (.A1(n_827_o_0),
    .A2(n_1361_o_0),
    .B(n_1362_o_0),
    .Y(n_1363_o_0));
 XNOR2xp5_ASAP7_75t_R n_1364 (.A(_00934_),
    .B(_00966_),
    .Y(n_1364_o_0));
 XOR2xp5_ASAP7_75t_R n_1365 (.A(_00424_),
    .B(_00870_),
    .Y(n_1365_o_0));
 NOR2xp33_ASAP7_75t_R n_1366 (.A(ld),
    .B(n_1365_o_0),
    .Y(n_1366_o_0));
 NAND2xp33_ASAP7_75t_R n_1367 (.A(_00902_),
    .B(n_1364_o_0),
    .Y(n_1367_o_0));
 OAI211xp5_ASAP7_75t_R n_1368 (.A1(_00902_),
    .A2(n_1364_o_0),
    .B(n_1366_o_0),
    .C(n_1367_o_0),
    .Y(n_1368_o_0));
 OAI21xp33_ASAP7_75t_R n_1369 (.A1(_00902_),
    .A2(n_1364_o_0),
    .B(n_1367_o_0),
    .Y(n_1369_o_0));
 AND2x2_ASAP7_75t_R n_1370 (.A(n_827_o_0),
    .B(n_1365_o_0),
    .Y(n_1370_o_0));
 AOI22xp33_ASAP7_75t_R n_1371 (.A1(n_1369_o_0),
    .A2(n_1370_o_0),
    .B1(key[10]),
    .B2(ld),
    .Y(n_1371_o_0));
 NAND2x1p5_ASAP7_75t_R n_1372 (.A(n_1371_o_0),
    .B(n_1368_o_0),
    .Y(n_1372_o_0));
 XNOR2xp5_ASAP7_75t_R n_1373 (.A(_00433_),
    .B(_00869_),
    .Y(n_1373_o_0));
 NAND2xp33_ASAP7_75t_R n_1374 (.A(_00901_),
    .B(n_1373_o_0),
    .Y(n_1374_o_0));
 OAI21xp33_ASAP7_75t_R n_1375 (.A1(_00901_),
    .A2(n_1373_o_0),
    .B(n_1374_o_0),
    .Y(n_1375_o_0));
 XNOR2xp5_ASAP7_75t_R n_1376 (.A(_00933_),
    .B(_00965_),
    .Y(n_1376_o_0));
 NAND2xp33_ASAP7_75t_R n_1377 (.A(n_1376_o_0),
    .B(n_1375_o_0),
    .Y(n_1377_o_0));
 OAI21xp33_ASAP7_75t_R n_1378 (.A1(n_1375_o_0),
    .A2(n_1376_o_0),
    .B(n_1377_o_0),
    .Y(n_1378_o_0));
 NAND2xp33_ASAP7_75t_R n_1379 (.A(key[9]),
    .B(ld),
    .Y(n_1379_o_0));
 OAI21xp5_ASAP7_75t_R n_1380 (.A1(ld),
    .A2(n_1378_o_0),
    .B(n_1379_o_0),
    .Y(n_1380_o_0));
 XNOR2xp5_ASAP7_75t_R n_1381 (.A(_00932_),
    .B(_00964_),
    .Y(n_1381_o_0));
 XNOR2xp5_ASAP7_75t_R n_1382 (.A(_00432_),
    .B(_00868_),
    .Y(n_1382_o_0));
 NAND2xp33_ASAP7_75t_R n_1383 (.A(_00900_),
    .B(n_1382_o_0),
    .Y(n_1383_o_0));
 OAI21xp33_ASAP7_75t_R n_1384 (.A1(_00900_),
    .A2(n_1382_o_0),
    .B(n_1383_o_0),
    .Y(n_1384_o_0));
 XNOR2xp5_ASAP7_75t_R n_1385 (.A(n_1381_o_0),
    .B(n_1384_o_0),
    .Y(n_1385_o_0));
 NOR2xp33_ASAP7_75t_R n_1386 (.A(key[8]),
    .B(n_827_o_0),
    .Y(n_1386_o_0));
 AOI21x1_ASAP7_75t_R n_1387 (.A1(n_827_o_0),
    .A2(n_1385_o_0),
    .B(n_1386_o_0),
    .Y(n_1387_o_0));
 NAND2xp33_ASAP7_75t_R n_1388 (.A(n_1380_o_0),
    .B(n_1387_o_0),
    .Y(n_1388_o_0));
 AO21x1_ASAP7_75t_R n_1389 (.A1(n_1385_o_0),
    .A2(n_827_o_0),
    .B(n_1386_o_0),
    .Y(n_1389_o_0));
 NOR2xp33_ASAP7_75t_R n_1390 (.A(n_1372_o_0),
    .B(n_1389_o_0),
    .Y(n_1390_o_0));
 XNOR2xp5_ASAP7_75t_R n_1391 (.A(_00935_),
    .B(_00967_),
    .Y(n_1391_o_0));
 XOR2xp5_ASAP7_75t_R n_1392 (.A(_00434_),
    .B(_00871_),
    .Y(n_1392_o_0));
 INVx1_ASAP7_75t_R n_1393 (.A(_00903_),
    .Y(n_1393_o_0));
 NAND2xp33_ASAP7_75t_R n_1394 (.A(n_1393_o_0),
    .B(n_1392_o_0),
    .Y(n_1394_o_0));
 OAI21xp33_ASAP7_75t_R n_1395 (.A1(n_1392_o_0),
    .A2(n_1393_o_0),
    .B(n_1394_o_0),
    .Y(n_1395_o_0));
 XNOR2xp5_ASAP7_75t_R n_1396 (.A(n_1391_o_0),
    .B(n_1395_o_0),
    .Y(n_1396_o_0));
 NOR2xp33_ASAP7_75t_R n_1397 (.A(key[11]),
    .B(n_827_o_0),
    .Y(n_1397_o_0));
 AOI21x1_ASAP7_75t_R n_1398 (.A1(n_827_o_0),
    .A2(n_1396_o_0),
    .B(n_1397_o_0),
    .Y(n_1398_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1399 (.A1(n_1372_o_0),
    .A2(n_1388_o_0),
    .B(n_1390_o_0),
    .C(n_1398_o_0),
    .Y(n_1399_o_0));
 NOR2xp33_ASAP7_75t_R n_1400 (.A(n_1363_o_0),
    .B(n_1399_o_0),
    .Y(n_1400_o_0));
 INVx1_ASAP7_75t_R n_1401 (.A(n_1400_o_0),
    .Y(n_1401_o_0));
 OR2x2_ASAP7_75t_R n_1402 (.A(n_1376_o_0),
    .B(n_1375_o_0),
    .Y(n_1402_o_0));
 INVx1_ASAP7_75t_R n_1403 (.A(n_1379_o_0),
    .Y(n_1403_o_0));
 AOI31xp67_ASAP7_75t_R n_1404 (.A1(n_827_o_0),
    .A2(n_1402_o_0),
    .A3(n_1377_o_0),
    .B(n_1403_o_0),
    .Y(n_1404_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1405 (.A1(n_827_o_0),
    .A2(n_1385_o_0),
    .B(n_1386_o_0),
    .C(n_1404_o_0),
    .Y(n_1405_o_0));
 OAI21xp33_ASAP7_75t_R n_1406 (.A1(n_1404_o_0),
    .A2(n_1389_o_0),
    .B(n_1405_o_0),
    .Y(n_1406_o_0));
 INVx1_ASAP7_75t_R n_1407 (.A(n_1398_o_0),
    .Y(n_1407_o_0));
 AOI21xp33_ASAP7_75t_R n_1408 (.A1(n_1372_o_0),
    .A2(n_1406_o_0),
    .B(n_1407_o_0),
    .Y(n_1408_o_0));
 NOR2xp33_ASAP7_75t_R n_1409 (.A(n_1380_o_0),
    .B(n_1389_o_0),
    .Y(n_1409_o_0));
 INVx1_ASAP7_75t_R n_1410 (.A(n_1409_o_0),
    .Y(n_1410_o_0));
 INVx1_ASAP7_75t_R n_1411 (.A(n_1372_o_0),
    .Y(n_1411_o_0));
 NOR3xp33_ASAP7_75t_R n_1412 (.A(n_1410_o_0),
    .B(net71),
    .C(net28),
    .Y(n_1412_o_0));
 OAI21xp33_ASAP7_75t_R n_1413 (.A1(n_1408_o_0),
    .A2(n_1412_o_0),
    .B(n_1363_o_0),
    .Y(n_1413_o_0));
 NAND2xp33_ASAP7_75t_R n_1414 (.A(n_1368_o_0),
    .B(n_1371_o_0),
    .Y(n_1414_o_0));
 INVx1_ASAP7_75t_R n_1415 (.A(n_1414_o_0),
    .Y(n_1415_o_0));
 NOR2xp33_ASAP7_75t_R n_1416 (.A(n_1387_o_0),
    .B(n_1404_o_0),
    .Y(n_1416_o_0));
 NAND2xp33_ASAP7_75t_R n_1417 (.A(n_1415_o_0),
    .B(n_1416_o_0),
    .Y(n_1417_o_0));
 INVx1_ASAP7_75t_R n_1418 (.A(n_1417_o_0),
    .Y(n_1418_o_0));
 XOR2xp5_ASAP7_75t_R n_1419 (.A(_00436_),
    .B(_00873_),
    .Y(n_1419_o_0));
 XNOR2xp5_ASAP7_75t_R n_1420 (.A(_00905_),
    .B(n_1419_o_0),
    .Y(n_1420_o_0));
 XNOR2xp5_ASAP7_75t_R n_1421 (.A(_00937_),
    .B(n_1420_o_0),
    .Y(n_1421_o_0));
 INVx1_ASAP7_75t_R n_1422 (.A(_00969_),
    .Y(n_1422_o_0));
 NAND2xp33_ASAP7_75t_R n_1423 (.A(n_1422_o_0),
    .B(n_1421_o_0),
    .Y(n_1423_o_0));
 OAI21xp33_ASAP7_75t_R n_1424 (.A1(n_1421_o_0),
    .A2(n_1422_o_0),
    .B(n_1423_o_0),
    .Y(n_1424_o_0));
 NAND2xp33_ASAP7_75t_R n_1425 (.A(key[13]),
    .B(ld),
    .Y(n_1425_o_0));
 OAI21xp5_ASAP7_75t_R n_1426 (.A1(ld),
    .A2(n_1424_o_0),
    .B(n_1425_o_0),
    .Y(n_1426_o_0));
 AOI21xp33_ASAP7_75t_R n_1427 (.A1(net13),
    .A2(n_1418_o_0),
    .B(n_1426_o_0),
    .Y(n_1427_o_0));
 NAND2xp33_ASAP7_75t_R n_1428 (.A(n_1372_o_0),
    .B(n_1387_o_0),
    .Y(n_1428_o_0));
 NAND2xp33_ASAP7_75t_R n_1429 (.A(n_1398_o_0),
    .B(n_1428_o_0),
    .Y(n_1429_o_0));
 AOI21xp33_ASAP7_75t_R n_1430 (.A1(n_1372_o_0),
    .A2(n_1404_o_0),
    .B(n_1398_o_0),
    .Y(n_1430_o_0));
 NAND2xp33_ASAP7_75t_R n_1431 (.A(n_1411_o_0),
    .B(n_1406_o_0),
    .Y(n_1431_o_0));
 AOI21xp33_ASAP7_75t_R n_1432 (.A1(n_1430_o_0),
    .A2(n_1431_o_0),
    .B(n_1363_o_0),
    .Y(n_1432_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1433 (.A1(net28),
    .A2(n_1410_o_0),
    .B(n_1429_o_0),
    .C(n_1432_o_0),
    .Y(n_1433_o_0));
 NAND2xp33_ASAP7_75t_R n_1434 (.A(n_1380_o_0),
    .B(n_1389_o_0),
    .Y(n_1434_o_0));
 AOI21xp33_ASAP7_75t_R n_1435 (.A1(net99),
    .A2(n_1434_o_0),
    .B(n_1407_o_0),
    .Y(n_1435_o_0));
 NOR2xp67_ASAP7_75t_R n_1436 (.A(n_1380_o_0),
    .B(n_1387_o_0),
    .Y(n_1436_o_0));
 NAND3xp33_ASAP7_75t_R n_1437 (.A(n_1436_o_0),
    .B(n_1407_o_0),
    .C(n_1372_o_0),
    .Y(n_1437_o_0));
 NOR2xp33_ASAP7_75t_R n_1438 (.A(n_1372_o_0),
    .B(n_1436_o_0),
    .Y(n_1438_o_0));
 INVx1_ASAP7_75t_R n_1439 (.A(n_1438_o_0),
    .Y(n_1439_o_0));
 AOI21xp33_ASAP7_75t_R n_1440 (.A1(n_1437_o_0),
    .A2(n_1439_o_0),
    .B(net71),
    .Y(n_1440_o_0));
 OAI21xp33_ASAP7_75t_R n_1441 (.A1(n_1435_o_0),
    .A2(n_1440_o_0),
    .B(n_1363_o_0),
    .Y(n_1441_o_0));
 AOI33xp33_ASAP7_75t_R n_1442 (.A1(n_1401_o_0),
    .A2(n_1413_o_0),
    .A3(n_1427_o_0),
    .B1(n_1433_o_0),
    .B2(n_1441_o_0),
    .B3(n_1426_o_0),
    .Y(n_1442_o_0));
 NOR2xp33_ASAP7_75t_R n_1443 (.A(ld),
    .B(n_1354_o_0),
    .Y(n_1443_o_0));
 NOR2xp33_ASAP7_75t_R n_1444 (.A(key[14]),
    .B(n_827_o_0),
    .Y(n_1444_o_0));
 INVx1_ASAP7_75t_R n_1445 (.A(n_1437_o_0),
    .Y(n_1445_o_0));
 OAI31xp33_ASAP7_75t_R n_1446 (.A1(n_1411_o_0),
    .A2(n_1404_o_0),
    .A3(n_1387_o_0),
    .B(n_1398_o_0),
    .Y(n_1446_o_0));
 OAI21xp33_ASAP7_75t_R n_1447 (.A1(n_1380_o_0),
    .A2(n_1389_o_0),
    .B(n_1411_o_0),
    .Y(n_1447_o_0));
 INVx1_ASAP7_75t_R n_1448 (.A(n_1447_o_0),
    .Y(n_1448_o_0));
 AO21x1_ASAP7_75t_R n_1449 (.A1(n_1361_o_0),
    .A2(n_827_o_0),
    .B(n_1362_o_0),
    .Y(n_1449_o_0));
 OAI21xp33_ASAP7_75t_R n_1450 (.A1(n_1446_o_0),
    .A2(n_1448_o_0),
    .B(n_1449_o_0),
    .Y(n_1450_o_0));
 NAND3xp33_ASAP7_75t_R n_1451 (.A(n_1410_o_0),
    .B(net44),
    .C(net28),
    .Y(n_1451_o_0));
 NOR2xp33_ASAP7_75t_R n_1452 (.A(n_1411_o_0),
    .B(n_1407_o_0),
    .Y(n_1452_o_0));
 NAND2xp33_ASAP7_75t_R n_1453 (.A(n_1436_o_0),
    .B(n_1452_o_0),
    .Y(n_1453_o_0));
 NOR3xp33_ASAP7_75t_R n_1454 (.A(n_1416_o_0),
    .B(n_1411_o_0),
    .C(n_1398_o_0),
    .Y(n_1454_o_0));
 INVx1_ASAP7_75t_R n_1455 (.A(n_1454_o_0),
    .Y(n_1455_o_0));
 NAND4xp25_ASAP7_75t_R n_1456 (.A(n_1451_o_0),
    .B(n_1453_o_0),
    .C(n_1455_o_0),
    .D(n_1363_o_0),
    .Y(n_1456_o_0));
 OAI211xp5_ASAP7_75t_R n_1457 (.A1(n_1445_o_0),
    .A2(n_1450_o_0),
    .B(n_1456_o_0),
    .C(n_1426_o_0),
    .Y(n_1457_o_0));
 NOR3xp33_ASAP7_75t_R n_1458 (.A(n_1436_o_0),
    .B(n_1407_o_0),
    .C(n_1411_o_0),
    .Y(n_1458_o_0));
 NOR2xp33_ASAP7_75t_R n_1459 (.A(n_1363_o_0),
    .B(n_1458_o_0),
    .Y(n_1459_o_0));
 OAI31xp33_ASAP7_75t_R n_1460 (.A1(n_1389_o_0),
    .A2(net99),
    .A3(net13),
    .B(n_1459_o_0),
    .Y(n_1460_o_0));
 NAND2xp33_ASAP7_75t_R n_1461 (.A(n_1372_o_0),
    .B(n_1416_o_0),
    .Y(n_1461_o_0));
 INVx1_ASAP7_75t_R n_1462 (.A(n_1461_o_0),
    .Y(n_1462_o_0));
 NAND2xp33_ASAP7_75t_R n_1463 (.A(n_1387_o_0),
    .B(n_1411_o_0),
    .Y(n_1463_o_0));
 INVx1_ASAP7_75t_R n_1464 (.A(n_1463_o_0),
    .Y(n_1464_o_0));
 NOR3xp33_ASAP7_75t_R n_1465 (.A(n_1462_o_0),
    .B(n_1464_o_0),
    .C(net71),
    .Y(n_1465_o_0));
 NAND2xp33_ASAP7_75t_R n_1466 (.A(n_1372_o_0),
    .B(n_1380_o_0),
    .Y(n_1466_o_0));
 NOR2xp33_ASAP7_75t_R n_1467 (.A(n_1414_o_0),
    .B(n_1406_o_0),
    .Y(n_1467_o_0));
 AOI21xp33_ASAP7_75t_R n_1468 (.A1(net13),
    .A2(n_1467_o_0),
    .B(n_1449_o_0),
    .Y(n_1468_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1469 (.A1(net20),
    .A2(n_1466_o_0),
    .B(n_1468_o_0),
    .C(n_1426_o_0),
    .Y(n_1469_o_0));
 OAI21xp33_ASAP7_75t_R n_1470 (.A1(n_1460_o_0),
    .A2(n_1465_o_0),
    .B(n_1469_o_0),
    .Y(n_1470_o_0));
 OAI211xp5_ASAP7_75t_R n_1471 (.A1(n_1443_o_0),
    .A2(n_1444_o_0),
    .B(n_1457_o_0),
    .C(n_1470_o_0),
    .Y(n_1471_o_0));
 OAI21xp33_ASAP7_75t_R n_1472 (.A1(n_1355_o_0),
    .A2(n_1442_o_0),
    .B(n_1471_o_0),
    .Y(n_1472_o_0));
 INVx1_ASAP7_75t_R n_1473 (.A(n_1436_o_0),
    .Y(n_1473_o_0));
 OAI21xp33_ASAP7_75t_R n_1474 (.A1(net99),
    .A2(n_1473_o_0),
    .B(n_1408_o_0),
    .Y(n_1474_o_0));
 OAI211xp5_ASAP7_75t_R n_1475 (.A1(n_1380_o_0),
    .A2(n_1387_o_0),
    .B(n_1407_o_0),
    .C(n_1372_o_0),
    .Y(n_1475_o_0));
 AND3x1_ASAP7_75t_R n_1476 (.A(n_1474_o_0),
    .B(n_1451_o_0),
    .C(n_1475_o_0),
    .Y(n_1476_o_0));
 NAND2xp33_ASAP7_75t_R n_1477 (.A(n_1380_o_0),
    .B(n_1387_o_0),
    .Y(n_1477_o_0));
 AOI31xp33_ASAP7_75t_R n_1478 (.A1(n_1405_o_0),
    .A2(n_1477_o_0),
    .A3(n_1372_o_0),
    .B(n_1398_o_0),
    .Y(n_1478_o_0));
 OAI21xp33_ASAP7_75t_R n_1479 (.A1(n_1404_o_0),
    .A2(net99),
    .B(n_1478_o_0),
    .Y(n_1479_o_0));
 NOR2xp33_ASAP7_75t_R n_1480 (.A(n_1380_o_0),
    .B(n_1387_o_0),
    .Y(n_1480_o_0));
 AOI211xp5_ASAP7_75t_R n_1481 (.A1(n_827_o_0),
    .A2(n_1385_o_0),
    .B(n_1404_o_0),
    .C(n_1386_o_0),
    .Y(n_1481_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1482 (.A1(n_1480_o_0),
    .A2(n_1481_o_0),
    .B(n_1411_o_0),
    .C(n_1407_o_0),
    .Y(n_1482_o_0));
 NOR3xp33_ASAP7_75t_R n_1483 (.A(n_1482_o_0),
    .B(n_1449_o_0),
    .C(n_1426_o_0),
    .Y(n_1483_o_0));
 INVx1_ASAP7_75t_R n_1484 (.A(n_1355_o_0),
    .Y(n_1484_o_0));
 AOI21xp33_ASAP7_75t_R n_1485 (.A1(n_1479_o_0),
    .A2(n_1483_o_0),
    .B(n_1484_o_0),
    .Y(n_1485_o_0));
 OAI31xp33_ASAP7_75t_R n_1486 (.A1(n_1426_o_0),
    .A2(n_1476_o_0),
    .A3(n_1363_o_0),
    .B(n_1485_o_0),
    .Y(n_1486_o_0));
 NOR2xp33_ASAP7_75t_R n_1487 (.A(n_1414_o_0),
    .B(n_1388_o_0),
    .Y(n_1487_o_0));
 INVx1_ASAP7_75t_R n_1488 (.A(n_1487_o_0),
    .Y(n_1488_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1489 (.A1(n_1480_o_0),
    .A2(n_1481_o_0),
    .B(n_1372_o_0),
    .C(n_1398_o_0),
    .Y(n_1489_o_0));
 AOI21xp33_ASAP7_75t_R n_1490 (.A1(net99),
    .A2(n_1410_o_0),
    .B(n_1438_o_0),
    .Y(n_1490_o_0));
 OAI21xp33_ASAP7_75t_R n_1491 (.A1(net13),
    .A2(n_1490_o_0),
    .B(n_1449_o_0),
    .Y(n_1491_o_0));
 AOI21xp33_ASAP7_75t_R n_1492 (.A1(n_1488_o_0),
    .A2(n_1489_o_0),
    .B(n_1491_o_0),
    .Y(n_1492_o_0));
 INVx1_ASAP7_75t_R n_1493 (.A(n_1421_o_0),
    .Y(n_1493_o_0));
 NAND2xp33_ASAP7_75t_R n_1494 (.A(_00969_),
    .B(n_1493_o_0),
    .Y(n_1494_o_0));
 INVx1_ASAP7_75t_R n_1495 (.A(n_1425_o_0),
    .Y(n_1495_o_0));
 AOI31xp67_ASAP7_75t_R n_1496 (.A1(n_827_o_0),
    .A2(n_1494_o_0),
    .A3(n_1423_o_0),
    .B(n_1495_o_0),
    .Y(n_1496_o_0));
 NAND2xp33_ASAP7_75t_R n_1497 (.A(n_1407_o_0),
    .B(n_1428_o_0),
    .Y(n_1497_o_0));
 INVx1_ASAP7_75t_R n_1498 (.A(n_1497_o_0),
    .Y(n_1498_o_0));
 NOR2xp33_ASAP7_75t_R n_1499 (.A(n_1380_o_0),
    .B(n_1387_o_0),
    .Y(n_1499_o_0));
 INVx1_ASAP7_75t_R n_1500 (.A(n_1499_o_0),
    .Y(n_1500_o_0));
 INVx1_ASAP7_75t_R n_1501 (.A(n_1428_o_0),
    .Y(n_1501_o_0));
 OAI21xp33_ASAP7_75t_R n_1502 (.A1(n_1499_o_0),
    .A2(n_1501_o_0),
    .B(n_1398_o_0),
    .Y(n_1502_o_0));
 INVx1_ASAP7_75t_R n_1503 (.A(n_1502_o_0),
    .Y(n_1503_o_0));
 AOI211xp5_ASAP7_75t_R n_1504 (.A1(n_1498_o_0),
    .A2(n_1500_o_0),
    .B(n_1503_o_0),
    .C(n_1449_o_0),
    .Y(n_1504_o_0));
 NOR3xp33_ASAP7_75t_R n_1505 (.A(n_1492_o_0),
    .B(n_1496_o_0),
    .C(n_1504_o_0),
    .Y(n_1505_o_0));
 AO21x1_ASAP7_75t_R n_1506 (.A1(n_1435_o_0),
    .A2(n_1417_o_0),
    .B(n_1363_o_0),
    .Y(n_1506_o_0));
 NOR2xp33_ASAP7_75t_R n_1507 (.A(n_1372_o_0),
    .B(n_1387_o_0),
    .Y(n_1507_o_0));
 NOR2xp33_ASAP7_75t_R n_1508 (.A(n_1398_o_0),
    .B(n_1507_o_0),
    .Y(n_1508_o_0));
 AOI21xp33_ASAP7_75t_R n_1509 (.A1(n_1372_o_0),
    .A2(n_1389_o_0),
    .B(n_1398_o_0),
    .Y(n_1509_o_0));
 INVx1_ASAP7_75t_R n_1510 (.A(n_1509_o_0),
    .Y(n_1510_o_0));
 NAND2xp33_ASAP7_75t_R n_1511 (.A(n_1411_o_0),
    .B(n_1388_o_0),
    .Y(n_1511_o_0));
 AOI21xp33_ASAP7_75t_R n_1512 (.A1(n_1511_o_0),
    .A2(n_1408_o_0),
    .B(n_1449_o_0),
    .Y(n_1512_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1513 (.A1(n_1418_o_0),
    .A2(n_1510_o_0),
    .B(n_1512_o_0),
    .C(n_1496_o_0),
    .Y(n_1513_o_0));
 OAI21xp33_ASAP7_75t_R n_1514 (.A1(n_1506_o_0),
    .A2(n_1508_o_0),
    .B(n_1513_o_0),
    .Y(n_1514_o_0));
 AOI21xp33_ASAP7_75t_R n_1515 (.A1(n_1380_o_0),
    .A2(n_1387_o_0),
    .B(n_1411_o_0),
    .Y(n_1515_o_0));
 OAI211xp5_ASAP7_75t_R n_1516 (.A1(n_1380_o_0),
    .A2(net28),
    .B(n_1417_o_0),
    .C(net44),
    .Y(n_1516_o_0));
 OAI31xp33_ASAP7_75t_R n_1517 (.A1(n_1507_o_0),
    .A2(n_1515_o_0),
    .A3(net20),
    .B(n_1516_o_0),
    .Y(n_1517_o_0));
 NAND3xp33_ASAP7_75t_R n_1518 (.A(n_1407_o_0),
    .B(n_1404_o_0),
    .C(n_1411_o_0),
    .Y(n_1518_o_0));
 NAND4xp25_ASAP7_75t_R n_1519 (.A(n_1399_o_0),
    .B(n_1518_o_0),
    .C(n_1437_o_0),
    .D(n_1449_o_0),
    .Y(n_1519_o_0));
 OAI211xp5_ASAP7_75t_R n_1520 (.A1(n_1517_o_0),
    .A2(n_1449_o_0),
    .B(n_1496_o_0),
    .C(n_1519_o_0),
    .Y(n_1520_o_0));
 INVx1_ASAP7_75t_R n_1521 (.A(n_1347_o_0),
    .Y(n_1521_o_0));
 AOI31xp33_ASAP7_75t_R n_1522 (.A1(n_1484_o_0),
    .A2(n_1514_o_0),
    .A3(n_1520_o_0),
    .B(n_1521_o_0),
    .Y(n_1522_o_0));
 OAI21xp33_ASAP7_75t_R n_1523 (.A1(n_1486_o_0),
    .A2(n_1505_o_0),
    .B(n_1522_o_0),
    .Y(n_1523_o_0));
 OAI21xp33_ASAP7_75t_R n_1524 (.A1(n_1347_o_0),
    .A2(n_1472_o_0),
    .B(n_1523_o_0),
    .Y(n_1524_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1525 (.A1(net28),
    .A2(n_1388_o_0),
    .B(n_1508_o_0),
    .C(n_1408_o_0),
    .Y(n_1525_o_0));
 OAI31xp33_ASAP7_75t_R n_1526 (.A1(n_1426_o_0),
    .A2(n_1525_o_0),
    .A3(n_1363_o_0),
    .B(n_1484_o_0),
    .Y(n_1526_o_0));
 OAI21xp33_ASAP7_75t_R n_1527 (.A1(n_1414_o_0),
    .A2(n_1436_o_0),
    .B(net44),
    .Y(n_1527_o_0));
 INVx1_ASAP7_75t_R n_1528 (.A(n_1406_o_0),
    .Y(n_1528_o_0));
 OAI21xp33_ASAP7_75t_R n_1529 (.A1(n_1414_o_0),
    .A2(n_1388_o_0),
    .B(n_1398_o_0),
    .Y(n_1529_o_0));
 AO21x1_ASAP7_75t_R n_1530 (.A1(n_1528_o_0),
    .A2(net99),
    .B(n_1529_o_0),
    .Y(n_1530_o_0));
 OA21x2_ASAP7_75t_R n_1531 (.A1(n_1527_o_0),
    .A2(n_1515_o_0),
    .B(n_1530_o_0),
    .Y(n_1531_o_0));
 AOI21xp33_ASAP7_75t_R n_1532 (.A1(n_1390_o_0),
    .A2(n_1407_o_0),
    .B(n_1496_o_0),
    .Y(n_1532_o_0));
 OAI31xp33_ASAP7_75t_R n_1533 (.A1(net20),
    .A2(n_1406_o_0),
    .A3(n_1414_o_0),
    .B(n_1532_o_0),
    .Y(n_1533_o_0));
 NOR3xp33_ASAP7_75t_R n_1534 (.A(n_1533_o_0),
    .B(n_1458_o_0),
    .C(n_1445_o_0),
    .Y(n_1534_o_0));
 AOI211xp5_ASAP7_75t_R n_1535 (.A1(n_1531_o_0),
    .A2(n_1496_o_0),
    .B(n_1534_o_0),
    .C(n_1449_o_0),
    .Y(n_1535_o_0));
 OAI21xp33_ASAP7_75t_R n_1536 (.A1(net99),
    .A2(n_1473_o_0),
    .B(n_1498_o_0),
    .Y(n_1536_o_0));
 OAI211xp5_ASAP7_75t_R n_1537 (.A1(n_1389_o_0),
    .A2(n_1411_o_0),
    .B(n_1398_o_0),
    .C(n_1380_o_0),
    .Y(n_1537_o_0));
 AOI211xp5_ASAP7_75t_R n_1538 (.A1(n_1536_o_0),
    .A2(n_1537_o_0),
    .B(n_1496_o_0),
    .C(n_1363_o_0),
    .Y(n_1538_o_0));
 NOR2xp33_ASAP7_75t_R n_1539 (.A(n_1372_o_0),
    .B(n_1380_o_0),
    .Y(n_1539_o_0));
 INVx1_ASAP7_75t_R n_1540 (.A(n_1539_o_0),
    .Y(n_1540_o_0));
 OAI31xp33_ASAP7_75t_R n_1541 (.A1(n_1414_o_0),
    .A2(n_1380_o_0),
    .A3(n_1389_o_0),
    .B(n_1407_o_0),
    .Y(n_1541_o_0));
 NOR2xp33_ASAP7_75t_R n_1542 (.A(n_1411_o_0),
    .B(n_1388_o_0),
    .Y(n_1542_o_0));
 NOR2xp33_ASAP7_75t_R n_1543 (.A(n_1541_o_0),
    .B(n_1542_o_0),
    .Y(n_1543_o_0));
 AOI31xp33_ASAP7_75t_R n_1544 (.A1(n_1496_o_0),
    .A2(n_1540_o_0),
    .A3(net71),
    .B(n_1543_o_0),
    .Y(n_1544_o_0));
 OAI21xp33_ASAP7_75t_R n_1545 (.A1(n_1414_o_0),
    .A2(n_1434_o_0),
    .B(n_1398_o_0),
    .Y(n_1545_o_0));
 OAI21xp33_ASAP7_75t_R n_1546 (.A1(n_1542_o_0),
    .A2(n_1545_o_0),
    .B(n_1426_o_0),
    .Y(n_1546_o_0));
 NOR2xp33_ASAP7_75t_R n_1547 (.A(n_1436_o_0),
    .B(n_1510_o_0),
    .Y(n_1547_o_0));
 OAI21xp33_ASAP7_75t_R n_1548 (.A1(n_1404_o_0),
    .A2(n_1372_o_0),
    .B(n_1498_o_0),
    .Y(n_1548_o_0));
 NAND3xp33_ASAP7_75t_R n_1549 (.A(n_1496_o_0),
    .B(n_1548_o_0),
    .C(n_1537_o_0),
    .Y(n_1549_o_0));
 OAI211xp5_ASAP7_75t_R n_1550 (.A1(n_1546_o_0),
    .A2(n_1547_o_0),
    .B(n_1549_o_0),
    .C(n_1363_o_0),
    .Y(n_1550_o_0));
 OAI21xp33_ASAP7_75t_R n_1551 (.A1(n_1363_o_0),
    .A2(n_1544_o_0),
    .B(n_1550_o_0),
    .Y(n_1551_o_0));
 OAI32xp33_ASAP7_75t_R n_1552 (.A1(n_1526_o_0),
    .A2(n_1535_o_0),
    .A3(n_1538_o_0),
    .B1(n_1551_o_0),
    .B2(n_1484_o_0),
    .Y(n_1552_o_0));
 AO21x1_ASAP7_75t_R n_1553 (.A1(n_1406_o_0),
    .A2(net28),
    .B(n_1515_o_0),
    .Y(n_1553_o_0));
 NOR2xp33_ASAP7_75t_R n_1554 (.A(net13),
    .B(n_1553_o_0),
    .Y(n_1554_o_0));
 NAND2xp33_ASAP7_75t_R n_1555 (.A(n_1372_o_0),
    .B(n_1404_o_0),
    .Y(n_1555_o_0));
 NAND2xp33_ASAP7_75t_R n_1556 (.A(n_1380_o_0),
    .B(n_1411_o_0),
    .Y(n_1556_o_0));
 OAI21xp33_ASAP7_75t_R n_1557 (.A1(net13),
    .A2(n_1556_o_0),
    .B(n_1363_o_0),
    .Y(n_1557_o_0));
 AOI21xp33_ASAP7_75t_R n_1558 (.A1(net20),
    .A2(n_1555_o_0),
    .B(n_1557_o_0),
    .Y(n_1558_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1559 (.A1(n_1454_o_0),
    .A2(n_1554_o_0),
    .B(n_1449_o_0),
    .C(n_1558_o_0),
    .Y(n_1559_o_0));
 NAND2xp33_ASAP7_75t_R n_1560 (.A(n_1426_o_0),
    .B(n_1449_o_0),
    .Y(n_1560_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1561 (.A1(n_1477_o_0),
    .A2(n_1405_o_0),
    .B(net28),
    .C(n_1398_o_0),
    .Y(n_1561_o_0));
 AOI21xp33_ASAP7_75t_R n_1562 (.A1(n_1372_o_0),
    .A2(n_1434_o_0),
    .B(n_1398_o_0),
    .Y(n_1562_o_0));
 AOI21xp33_ASAP7_75t_R n_1563 (.A1(n_1463_o_0),
    .A2(n_1562_o_0),
    .B(n_1496_o_0),
    .Y(n_1563_o_0));
 OAI21xp33_ASAP7_75t_R n_1564 (.A1(n_1561_o_0),
    .A2(n_1507_o_0),
    .B(n_1563_o_0),
    .Y(n_1564_o_0));
 NOR2xp33_ASAP7_75t_R n_1565 (.A(n_1414_o_0),
    .B(n_1416_o_0),
    .Y(n_1565_o_0));
 INVx1_ASAP7_75t_R n_1566 (.A(n_1565_o_0),
    .Y(n_1566_o_0));
 INVx1_ASAP7_75t_R n_1567 (.A(n_1466_o_0),
    .Y(n_1567_o_0));
 NOR3xp33_ASAP7_75t_R n_1568 (.A(n_1567_o_0),
    .B(n_1499_o_0),
    .C(net71),
    .Y(n_1568_o_0));
 INVx1_ASAP7_75t_R n_1569 (.A(n_1568_o_0),
    .Y(n_1569_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1570 (.A1(net20),
    .A2(n_1566_o_0),
    .B(n_1569_o_0),
    .C(n_1363_o_0),
    .Y(n_1570_o_0));
 AOI21xp33_ASAP7_75t_R n_1571 (.A1(n_1560_o_0),
    .A2(n_1564_o_0),
    .B(n_1570_o_0),
    .Y(n_1571_o_0));
 AOI21xp33_ASAP7_75t_R n_1572 (.A1(n_1427_o_0),
    .A2(n_1559_o_0),
    .B(n_1571_o_0),
    .Y(n_1572_o_0));
 NAND2xp33_ASAP7_75t_R n_1573 (.A(n_1407_o_0),
    .B(n_1463_o_0),
    .Y(n_1573_o_0));
 NOR2xp33_ASAP7_75t_R n_1574 (.A(net28),
    .B(n_1436_o_0),
    .Y(n_1574_o_0));
 AOI21xp33_ASAP7_75t_R n_1575 (.A1(n_1417_o_0),
    .A2(n_1408_o_0),
    .B(n_1449_o_0),
    .Y(n_1575_o_0));
 OAI21xp33_ASAP7_75t_R n_1576 (.A1(n_1387_o_0),
    .A2(n_1411_o_0),
    .B(n_1477_o_0),
    .Y(n_1576_o_0));
 AOI21xp33_ASAP7_75t_R n_1577 (.A1(net71),
    .A2(n_1576_o_0),
    .B(n_1509_o_0),
    .Y(n_1577_o_0));
 AOI211xp5_ASAP7_75t_R n_1578 (.A1(n_1467_o_0),
    .A2(net13),
    .B(n_1363_o_0),
    .C(n_1577_o_0),
    .Y(n_1578_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1579 (.A1(n_1573_o_0),
    .A2(n_1574_o_0),
    .B(n_1575_o_0),
    .C(n_1578_o_0),
    .Y(n_1579_o_0));
 OAI31xp33_ASAP7_75t_R n_1580 (.A1(n_1434_o_0),
    .A2(net28),
    .A3(net71),
    .B(n_1530_o_0),
    .Y(n_1580_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1581 (.A1(n_1387_o_0),
    .A2(n_1380_o_0),
    .B(n_1372_o_0),
    .C(n_1398_o_0),
    .Y(n_1581_o_0));
 AOI21xp33_ASAP7_75t_R n_1582 (.A1(n_1404_o_0),
    .A2(net99),
    .B(n_1581_o_0),
    .Y(n_1582_o_0));
 AOI31xp33_ASAP7_75t_R n_1583 (.A1(net99),
    .A2(net70),
    .A3(n_1388_o_0),
    .B(n_1582_o_0),
    .Y(n_1583_o_0));
 AOI31xp33_ASAP7_75t_R n_1584 (.A1(n_1426_o_0),
    .A2(n_1583_o_0),
    .A3(n_1363_o_0),
    .B(n_1355_o_0),
    .Y(n_1584_o_0));
 OAI21xp33_ASAP7_75t_R n_1585 (.A1(n_1560_o_0),
    .A2(n_1580_o_0),
    .B(n_1584_o_0),
    .Y(n_1585_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1586 (.A1(n_1496_o_0),
    .A2(n_1579_o_0),
    .B(n_1585_o_0),
    .C(n_1521_o_0),
    .Y(n_1586_o_0));
 AOI21xp33_ASAP7_75t_R n_1587 (.A1(n_1572_o_0),
    .A2(n_1355_o_0),
    .B(n_1586_o_0),
    .Y(n_1587_o_0));
 AOI21xp33_ASAP7_75t_R n_1588 (.A1(n_1347_o_0),
    .A2(n_1552_o_0),
    .B(n_1587_o_0),
    .Y(n_1588_o_0));
 NAND2xp33_ASAP7_75t_R n_1589 (.A(n_1407_o_0),
    .B(n_1417_o_0),
    .Y(n_1589_o_0));
 OAI21xp33_ASAP7_75t_R n_1590 (.A1(n_1567_o_0),
    .A2(net70),
    .B(n_1589_o_0),
    .Y(n_1590_o_0));
 AOI21xp33_ASAP7_75t_R n_1591 (.A1(n_1415_o_0),
    .A2(n_1416_o_0),
    .B(n_1407_o_0),
    .Y(n_1591_o_0));
 AOI21xp33_ASAP7_75t_R n_1592 (.A1(n_1591_o_0),
    .A2(n_1466_o_0),
    .B(n_1449_o_0),
    .Y(n_1592_o_0));
 OAI21xp33_ASAP7_75t_R n_1593 (.A1(n_1556_o_0),
    .A2(net71),
    .B(n_1592_o_0),
    .Y(n_1593_o_0));
 OAI21xp33_ASAP7_75t_R n_1594 (.A1(n_1363_o_0),
    .A2(n_1590_o_0),
    .B(n_1593_o_0),
    .Y(n_1594_o_0));
 OAI21xp33_ASAP7_75t_R n_1595 (.A1(n_1501_o_0),
    .A2(n_1529_o_0),
    .B(n_1363_o_0),
    .Y(n_1595_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1596 (.A1(n_1416_o_0),
    .A2(net99),
    .B(n_1408_o_0),
    .C(n_1363_o_0),
    .Y(n_1596_o_0));
 OAI31xp33_ASAP7_75t_R n_1597 (.A1(net28),
    .A2(net71),
    .A3(n_1436_o_0),
    .B(n_1596_o_0),
    .Y(n_1597_o_0));
 OAI211xp5_ASAP7_75t_R n_1598 (.A1(n_1543_o_0),
    .A2(n_1595_o_0),
    .B(n_1597_o_0),
    .C(n_1426_o_0),
    .Y(n_1598_o_0));
 OAI21xp33_ASAP7_75t_R n_1599 (.A1(n_1426_o_0),
    .A2(n_1594_o_0),
    .B(n_1598_o_0),
    .Y(n_1599_o_0));
 NOR3xp33_ASAP7_75t_R n_1600 (.A(n_1567_o_0),
    .B(n_1407_o_0),
    .C(n_1499_o_0),
    .Y(n_1600_o_0));
 INVx1_ASAP7_75t_R n_1601 (.A(n_1600_o_0),
    .Y(n_1601_o_0));
 OAI21xp33_ASAP7_75t_R n_1602 (.A1(net71),
    .A2(n_1539_o_0),
    .B(n_1601_o_0),
    .Y(n_1602_o_0));
 OAI31xp33_ASAP7_75t_R n_1603 (.A1(n_1480_o_0),
    .A2(n_1481_o_0),
    .A3(n_1414_o_0),
    .B(n_1398_o_0),
    .Y(n_1603_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1604 (.A1(n_1410_o_0),
    .A2(net99),
    .B(n_1603_o_0),
    .C(n_1363_o_0),
    .Y(n_1604_o_0));
 AOI31xp33_ASAP7_75t_R n_1605 (.A1(net20),
    .A2(n_1439_o_0),
    .A3(n_1466_o_0),
    .B(n_1604_o_0),
    .Y(n_1605_o_0));
 AOI21xp33_ASAP7_75t_R n_1606 (.A1(n_1449_o_0),
    .A2(n_1602_o_0),
    .B(n_1605_o_0),
    .Y(n_1606_o_0));
 AOI31xp33_ASAP7_75t_R n_1607 (.A1(n_1477_o_0),
    .A2(n_1405_o_0),
    .A3(n_1415_o_0),
    .B(n_1567_o_0),
    .Y(n_1607_o_0));
 AOI21xp33_ASAP7_75t_R n_1608 (.A1(n_1428_o_0),
    .A2(n_1556_o_0),
    .B(net44),
    .Y(n_1608_o_0));
 AO21x1_ASAP7_75t_R n_1609 (.A1(n_1607_o_0),
    .A2(net13),
    .B(n_1608_o_0),
    .Y(n_1609_o_0));
 AOI22xp33_ASAP7_75t_R n_1610 (.A1(n_1482_o_0),
    .A2(n_1461_o_0),
    .B1(net44),
    .B2(n_1567_o_0),
    .Y(n_1610_o_0));
 OAI21xp33_ASAP7_75t_R n_1611 (.A1(n_1363_o_0),
    .A2(n_1610_o_0),
    .B(n_1426_o_0),
    .Y(n_1611_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1612 (.A1(n_1363_o_0),
    .A2(n_1609_o_0),
    .B(n_1611_o_0),
    .C(n_1484_o_0),
    .Y(n_1612_o_0));
 AOI21xp33_ASAP7_75t_R n_1613 (.A1(n_1496_o_0),
    .A2(n_1606_o_0),
    .B(n_1612_o_0),
    .Y(n_1613_o_0));
 AOI21xp33_ASAP7_75t_R n_1614 (.A1(n_1355_o_0),
    .A2(n_1599_o_0),
    .B(n_1613_o_0),
    .Y(n_1614_o_0));
 AOI21xp33_ASAP7_75t_R n_1615 (.A1(n_1434_o_0),
    .A2(net99),
    .B(n_1545_o_0),
    .Y(n_1615_o_0));
 AOI21xp33_ASAP7_75t_R n_1616 (.A1(n_1607_o_0),
    .A2(net20),
    .B(n_1615_o_0),
    .Y(n_1616_o_0));
 AOI22xp33_ASAP7_75t_R n_1617 (.A1(n_1562_o_0),
    .A2(n_1511_o_0),
    .B1(n_1466_o_0),
    .B2(n_1591_o_0),
    .Y(n_1617_o_0));
 NAND3xp33_ASAP7_75t_R n_1618 (.A(n_1617_o_0),
    .B(n_1496_o_0),
    .C(n_1363_o_0),
    .Y(n_1618_o_0));
 OAI31xp33_ASAP7_75t_R n_1619 (.A1(n_1426_o_0),
    .A2(n_1616_o_0),
    .A3(n_1363_o_0),
    .B(n_1618_o_0),
    .Y(n_1619_o_0));
 OAI21xp33_ASAP7_75t_R n_1620 (.A1(n_1515_o_0),
    .A2(n_1529_o_0),
    .B(n_1589_o_0),
    .Y(n_1620_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1621 (.A1(n_1436_o_0),
    .A2(n_1415_o_0),
    .B(n_1429_o_0),
    .C(n_1363_o_0),
    .Y(n_1621_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1622 (.A1(n_1478_o_0),
    .A2(n_1540_o_0),
    .B(n_1621_o_0),
    .C(n_1426_o_0),
    .Y(n_1622_o_0));
 AOI21xp33_ASAP7_75t_R n_1623 (.A1(n_1620_o_0),
    .A2(n_1449_o_0),
    .B(n_1622_o_0),
    .Y(n_1623_o_0));
 NOR3xp33_ASAP7_75t_R n_1624 (.A(n_1619_o_0),
    .B(n_1623_o_0),
    .C(n_1484_o_0),
    .Y(n_1624_o_0));
 OAI21xp33_ASAP7_75t_R n_1625 (.A1(net99),
    .A2(n_1389_o_0),
    .B(n_1380_o_0),
    .Y(n_1625_o_0));
 NAND3xp33_ASAP7_75t_R n_1626 (.A(n_1416_o_0),
    .B(n_1407_o_0),
    .C(n_1415_o_0),
    .Y(n_1626_o_0));
 OAI21xp33_ASAP7_75t_R n_1627 (.A1(net13),
    .A2(n_1625_o_0),
    .B(n_1626_o_0),
    .Y(n_1627_o_0));
 INVx1_ASAP7_75t_R n_1628 (.A(n_1429_o_0),
    .Y(n_1628_o_0));
 OAI21xp33_ASAP7_75t_R n_1629 (.A1(n_1372_o_0),
    .A2(n_1388_o_0),
    .B(n_1407_o_0),
    .Y(n_1629_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1630 (.A1(n_1372_o_0),
    .A2(n_1409_o_0),
    .B(n_1629_o_0),
    .C(n_1363_o_0),
    .Y(n_1630_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1631 (.A1(n_1417_o_0),
    .A2(n_1628_o_0),
    .B(n_1630_o_0),
    .C(n_1496_o_0),
    .Y(n_1631_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1632 (.A1(n_1627_o_0),
    .A2(n_1412_o_0),
    .B(n_1449_o_0),
    .C(n_1631_o_0),
    .Y(n_1632_o_0));
 OAI22xp33_ASAP7_75t_R n_1633 (.A1(n_1467_o_0),
    .A2(n_1561_o_0),
    .B1(n_1510_o_0),
    .B2(n_1448_o_0),
    .Y(n_1633_o_0));
 AOI21xp33_ASAP7_75t_R n_1634 (.A1(n_1380_o_0),
    .A2(n_1387_o_0),
    .B(n_1497_o_0),
    .Y(n_1634_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1635 (.A1(n_1387_o_0),
    .A2(net28),
    .B(n_1404_o_0),
    .C(net44),
    .Y(n_1635_o_0));
 OAI31xp33_ASAP7_75t_R n_1636 (.A1(n_1449_o_0),
    .A2(n_1634_o_0),
    .A3(n_1635_o_0),
    .B(n_1426_o_0),
    .Y(n_1636_o_0));
 AOI21xp33_ASAP7_75t_R n_1637 (.A1(n_1633_o_0),
    .A2(n_1449_o_0),
    .B(n_1636_o_0),
    .Y(n_1637_o_0));
 NOR4xp25_ASAP7_75t_R n_1638 (.A(n_1632_o_0),
    .B(n_1637_o_0),
    .C(n_1355_o_0),
    .D(n_1521_o_0),
    .Y(n_1638_o_0));
 AOI21xp33_ASAP7_75t_R n_1639 (.A1(n_1347_o_0),
    .A2(n_1624_o_0),
    .B(n_1638_o_0),
    .Y(n_1639_o_0));
 OAI21xp33_ASAP7_75t_R n_1640 (.A1(n_1347_o_0),
    .A2(n_1614_o_0),
    .B(n_1639_o_0),
    .Y(n_1640_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1641 (.A1(n_1628_o_0),
    .A2(n_1447_o_0),
    .B(n_1543_o_0),
    .C(n_1449_o_0),
    .Y(n_1641_o_0));
 OAI211xp5_ASAP7_75t_R n_1642 (.A1(n_1449_o_0),
    .A2(n_1634_o_0),
    .B(n_1641_o_0),
    .C(n_1496_o_0),
    .Y(n_1642_o_0));
 INVx1_ASAP7_75t_R n_1643 (.A(n_1489_o_0),
    .Y(n_1643_o_0));
 INVx1_ASAP7_75t_R n_1644 (.A(n_1511_o_0),
    .Y(n_1644_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1645 (.A1(n_1409_o_0),
    .A2(n_1372_o_0),
    .B(n_1507_o_0),
    .C(n_1398_o_0),
    .Y(n_1645_o_0));
 OAI211xp5_ASAP7_75t_R n_1646 (.A1(n_1643_o_0),
    .A2(n_1644_o_0),
    .B(n_1645_o_0),
    .C(n_1363_o_0),
    .Y(n_1646_o_0));
 OAI21xp33_ASAP7_75t_R n_1647 (.A1(n_1568_o_0),
    .A2(n_1460_o_0),
    .B(n_1646_o_0),
    .Y(n_1647_o_0));
 AOI21xp33_ASAP7_75t_R n_1648 (.A1(n_1426_o_0),
    .A2(n_1647_o_0),
    .B(n_1355_o_0),
    .Y(n_1648_o_0));
 NAND2xp33_ASAP7_75t_R n_1649 (.A(n_1409_o_0),
    .B(n_1452_o_0),
    .Y(n_1649_o_0));
 NAND2xp33_ASAP7_75t_R n_1650 (.A(n_1426_o_0),
    .B(n_1649_o_0),
    .Y(n_1650_o_0));
 OAI21xp33_ASAP7_75t_R n_1651 (.A1(n_1387_o_0),
    .A2(net99),
    .B(n_1489_o_0),
    .Y(n_1651_o_0));
 OAI311xp33_ASAP7_75t_R n_1652 (.A1(net70),
    .A2(n_1644_o_0),
    .A3(n_1501_o_0),
    .B1(n_1496_o_0),
    .C1(n_1651_o_0),
    .Y(n_1652_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1653 (.A1(n_1447_o_0),
    .A2(n_1509_o_0),
    .B(n_1650_o_0),
    .C(n_1652_o_0),
    .Y(n_1653_o_0));
 NAND3xp33_ASAP7_75t_R n_1654 (.A(n_1406_o_0),
    .B(n_1407_o_0),
    .C(net99),
    .Y(n_1654_o_0));
 INVx1_ASAP7_75t_R n_1655 (.A(n_1654_o_0),
    .Y(n_1655_o_0));
 NAND2xp33_ASAP7_75t_R n_1656 (.A(n_1411_o_0),
    .B(n_1398_o_0),
    .Y(n_1656_o_0));
 AOI31xp33_ASAP7_75t_R n_1657 (.A1(n_1415_o_0),
    .A2(n_1404_o_0),
    .A3(n_1387_o_0),
    .B(n_1398_o_0),
    .Y(n_1657_o_0));
 AOI21xp33_ASAP7_75t_R n_1658 (.A1(n_1466_o_0),
    .A2(n_1657_o_0),
    .B(n_1426_o_0),
    .Y(n_1658_o_0));
 OAI21xp33_ASAP7_75t_R n_1659 (.A1(n_1656_o_0),
    .A2(n_1528_o_0),
    .B(n_1658_o_0),
    .Y(n_1659_o_0));
 OAI21xp33_ASAP7_75t_R n_1660 (.A1(n_1655_o_0),
    .A2(n_1496_o_0),
    .B(n_1659_o_0),
    .Y(n_1660_o_0));
 INVx1_ASAP7_75t_R n_1661 (.A(n_1656_o_0),
    .Y(n_1661_o_0));
 OAI21xp33_ASAP7_75t_R n_1662 (.A1(n_1567_o_0),
    .A2(n_1541_o_0),
    .B(n_1496_o_0),
    .Y(n_1662_o_0));
 AOI21xp33_ASAP7_75t_R n_1663 (.A1(n_1661_o_0),
    .A2(n_1406_o_0),
    .B(n_1662_o_0),
    .Y(n_1663_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1664 (.A1(n_1436_o_0),
    .A2(n_1452_o_0),
    .B(n_1449_o_0),
    .C(n_1355_o_0),
    .Y(n_1664_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1665 (.A1(n_1426_o_0),
    .A2(n_1654_o_0),
    .B(n_1663_o_0),
    .C(n_1664_o_0),
    .Y(n_1665_o_0));
 OAI21xp33_ASAP7_75t_R n_1666 (.A1(n_1355_o_0),
    .A2(n_1660_o_0),
    .B(n_1665_o_0),
    .Y(n_1666_o_0));
 AOI21xp33_ASAP7_75t_R n_1667 (.A1(n_1449_o_0),
    .A2(n_1653_o_0),
    .B(n_1666_o_0),
    .Y(n_1667_o_0));
 AOI21xp33_ASAP7_75t_R n_1668 (.A1(n_1642_o_0),
    .A2(n_1648_o_0),
    .B(n_1667_o_0),
    .Y(n_1668_o_0));
 NOR2xp33_ASAP7_75t_R n_1669 (.A(n_1372_o_0),
    .B(n_1416_o_0),
    .Y(n_1669_o_0));
 NAND2xp33_ASAP7_75t_R n_1670 (.A(n_1540_o_0),
    .B(n_1478_o_0),
    .Y(n_1670_o_0));
 OAI31xp33_ASAP7_75t_R n_1671 (.A1(n_1515_o_0),
    .A2(n_1669_o_0),
    .A3(net20),
    .B(n_1670_o_0),
    .Y(n_1671_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1672 (.A1(n_1410_o_0),
    .A2(net99),
    .B(n_1573_o_0),
    .C(n_1363_o_0),
    .Y(n_1672_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1673 (.A1(net28),
    .A2(n_1436_o_0),
    .B(n_1482_o_0),
    .C(n_1672_o_0),
    .Y(n_1673_o_0));
 AOI21xp33_ASAP7_75t_R n_1674 (.A1(n_1449_o_0),
    .A2(n_1671_o_0),
    .B(n_1673_o_0),
    .Y(n_1674_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1675 (.A1(n_1389_o_0),
    .A2(net99),
    .B(n_1404_o_0),
    .C(n_1405_o_0),
    .Y(n_1675_o_0));
 OAI211xp5_ASAP7_75t_R n_1676 (.A1(net71),
    .A2(n_1675_o_0),
    .B(n_1502_o_0),
    .C(n_1363_o_0),
    .Y(n_1676_o_0));
 OAI221xp5_ASAP7_75t_R n_1677 (.A1(n_1404_o_0),
    .A2(n_1389_o_0),
    .B1(n_1372_o_0),
    .B2(n_1405_o_0),
    .C(n_1407_o_0),
    .Y(n_1677_o_0));
 OAI31xp33_ASAP7_75t_R n_1678 (.A1(net28),
    .A2(n_1409_o_0),
    .A3(net70),
    .B(n_1677_o_0),
    .Y(n_1678_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1679 (.A1(n_1565_o_0),
    .A2(net71),
    .B(n_1678_o_0),
    .C(n_1449_o_0),
    .Y(n_1679_o_0));
 AO21x1_ASAP7_75t_R n_1680 (.A1(n_1676_o_0),
    .A2(n_1679_o_0),
    .B(n_1355_o_0),
    .Y(n_1680_o_0));
 OAI21xp33_ASAP7_75t_R n_1681 (.A1(n_1484_o_0),
    .A2(n_1674_o_0),
    .B(n_1680_o_0),
    .Y(n_1681_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1682 (.A1(n_1499_o_0),
    .A2(n_1464_o_0),
    .B(net44),
    .C(n_1363_o_0),
    .Y(n_1682_o_0));
 INVx1_ASAP7_75t_R n_1683 (.A(n_1682_o_0),
    .Y(n_1683_o_0));
 AOI21xp33_ASAP7_75t_R n_1684 (.A1(n_1447_o_0),
    .A2(n_1478_o_0),
    .B(n_1449_o_0),
    .Y(n_1684_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1685 (.A1(n_1404_o_0),
    .A2(net99),
    .B(n_1581_o_0),
    .C(n_1684_o_0),
    .Y(n_1685_o_0));
 OAI211xp5_ASAP7_75t_R n_1686 (.A1(n_1591_o_0),
    .A2(n_1683_o_0),
    .B(n_1685_o_0),
    .C(n_1484_o_0),
    .Y(n_1686_o_0));
 NAND2xp33_ASAP7_75t_R n_1687 (.A(n_1428_o_0),
    .B(n_1556_o_0),
    .Y(n_1687_o_0));
 AOI211xp5_ASAP7_75t_R n_1688 (.A1(net70),
    .A2(n_1687_o_0),
    .B(n_1482_o_0),
    .C(n_1449_o_0),
    .Y(n_1688_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1689 (.A1(n_1561_o_0),
    .A2(n_1539_o_0),
    .B(n_1682_o_0),
    .C(n_1688_o_0),
    .Y(n_1689_o_0));
 NAND2xp33_ASAP7_75t_R n_1690 (.A(n_1355_o_0),
    .B(n_1689_o_0),
    .Y(n_1690_o_0));
 AOI31xp33_ASAP7_75t_R n_1691 (.A1(n_1686_o_0),
    .A2(n_1690_o_0),
    .A3(n_1496_o_0),
    .B(n_1347_o_0),
    .Y(n_1691_o_0));
 OAI21xp33_ASAP7_75t_R n_1692 (.A1(n_1496_o_0),
    .A2(n_1681_o_0),
    .B(n_1691_o_0),
    .Y(n_1692_o_0));
 OAI21xp33_ASAP7_75t_R n_1693 (.A1(n_1521_o_0),
    .A2(n_1668_o_0),
    .B(n_1692_o_0),
    .Y(n_1693_o_0));
 AOI21xp33_ASAP7_75t_R n_1694 (.A1(n_1428_o_0),
    .A2(n_1540_o_0),
    .B(net20),
    .Y(n_1694_o_0));
 OAI21xp33_ASAP7_75t_R n_1695 (.A1(n_1694_o_0),
    .A2(n_1547_o_0),
    .B(n_1449_o_0),
    .Y(n_1695_o_0));
 OAI22xp33_ASAP7_75t_R n_1696 (.A1(n_1448_o_0),
    .A2(net20),
    .B1(n_1473_o_0),
    .B2(net28),
    .Y(n_1696_o_0));
 AOI21xp33_ASAP7_75t_R n_1697 (.A1(n_1363_o_0),
    .A2(n_1696_o_0),
    .B(n_1496_o_0),
    .Y(n_1697_o_0));
 AOI21xp33_ASAP7_75t_R n_1698 (.A1(n_1548_o_0),
    .A2(n_1601_o_0),
    .B(n_1363_o_0),
    .Y(n_1698_o_0));
 NAND2xp33_ASAP7_75t_R n_1699 (.A(n_1555_o_0),
    .B(n_1477_o_0),
    .Y(n_1699_o_0));
 OAI31xp33_ASAP7_75t_R n_1700 (.A1(net13),
    .A2(n_1438_o_0),
    .A3(n_1567_o_0),
    .B(n_1363_o_0),
    .Y(n_1700_o_0));
 AOI21xp33_ASAP7_75t_R n_1701 (.A1(net20),
    .A2(n_1699_o_0),
    .B(n_1700_o_0),
    .Y(n_1701_o_0));
 OAI31xp33_ASAP7_75t_R n_1702 (.A1(n_1698_o_0),
    .A2(n_1701_o_0),
    .A3(n_1426_o_0),
    .B(n_1484_o_0),
    .Y(n_1702_o_0));
 OAI31xp33_ASAP7_75t_R n_1703 (.A1(net13),
    .A2(n_1406_o_0),
    .A3(n_1414_o_0),
    .B(n_1626_o_0),
    .Y(n_1703_o_0));
 AOI211xp5_ASAP7_75t_R n_1704 (.A1(net99),
    .A2(n_1409_o_0),
    .B(n_1703_o_0),
    .C(n_1449_o_0),
    .Y(n_1704_o_0));
 NOR2xp33_ASAP7_75t_R n_1705 (.A(n_1398_o_0),
    .B(n_1515_o_0),
    .Y(n_1705_o_0));
 AOI21xp33_ASAP7_75t_R n_1706 (.A1(n_1705_o_0),
    .A2(n_1431_o_0),
    .B(n_1450_o_0),
    .Y(n_1706_o_0));
 NAND2xp33_ASAP7_75t_R n_1707 (.A(n_1511_o_0),
    .B(n_1562_o_0),
    .Y(n_1707_o_0));
 OAI31xp33_ASAP7_75t_R n_1708 (.A1(n_1462_o_0),
    .A2(n_1539_o_0),
    .A3(net13),
    .B(n_1707_o_0),
    .Y(n_1708_o_0));
 NAND3xp33_ASAP7_75t_R n_1709 (.A(n_1398_o_0),
    .B(n_1411_o_0),
    .C(n_1380_o_0),
    .Y(n_1709_o_0));
 NAND3xp33_ASAP7_75t_R n_1710 (.A(n_1455_o_0),
    .B(n_1709_o_0),
    .C(n_1626_o_0),
    .Y(n_1710_o_0));
 INVx1_ASAP7_75t_R n_1711 (.A(n_1459_o_0),
    .Y(n_1711_o_0));
 OAI221xp5_ASAP7_75t_R n_1712 (.A1(n_1449_o_0),
    .A2(n_1708_o_0),
    .B1(n_1710_o_0),
    .B2(n_1711_o_0),
    .C(n_1496_o_0),
    .Y(n_1712_o_0));
 OAI31xp33_ASAP7_75t_R n_1713 (.A1(n_1704_o_0),
    .A2(n_1706_o_0),
    .A3(n_1496_o_0),
    .B(n_1712_o_0),
    .Y(n_1713_o_0));
 AOI21xp33_ASAP7_75t_R n_1714 (.A1(n_1355_o_0),
    .A2(n_1713_o_0),
    .B(n_1347_o_0),
    .Y(n_1714_o_0));
 OAI21xp33_ASAP7_75t_R n_1715 (.A1(net13),
    .A2(n_1467_o_0),
    .B(n_1449_o_0),
    .Y(n_1715_o_0));
 AOI21xp33_ASAP7_75t_R n_1716 (.A1(net13),
    .A2(n_1388_o_0),
    .B(n_1715_o_0),
    .Y(n_1716_o_0));
 OAI211xp5_ASAP7_75t_R n_1717 (.A1(n_1380_o_0),
    .A2(n_1411_o_0),
    .B(n_1447_o_0),
    .C(n_1398_o_0),
    .Y(n_1717_o_0));
 AND3x1_ASAP7_75t_R n_1718 (.A(n_1455_o_0),
    .B(n_1717_o_0),
    .C(n_1363_o_0),
    .Y(n_1718_o_0));
 AOI21xp33_ASAP7_75t_R n_1719 (.A1(net13),
    .A2(n_1699_o_0),
    .B(n_1449_o_0),
    .Y(n_1719_o_0));
 OAI21xp33_ASAP7_75t_R n_1720 (.A1(n_1429_o_0),
    .A2(n_1448_o_0),
    .B(n_1719_o_0),
    .Y(n_1720_o_0));
 OAI311xp33_ASAP7_75t_R n_1721 (.A1(n_1503_o_0),
    .A2(n_1440_o_0),
    .A3(n_1363_o_0),
    .B1(n_1720_o_0),
    .C1(n_1496_o_0),
    .Y(n_1721_o_0));
 OAI31xp33_ASAP7_75t_R n_1722 (.A1(n_1716_o_0),
    .A2(n_1718_o_0),
    .A3(n_1496_o_0),
    .B(n_1721_o_0),
    .Y(n_1722_o_0));
 NOR2xp33_ASAP7_75t_R n_1723 (.A(n_1363_o_0),
    .B(n_1426_o_0),
    .Y(n_1723_o_0));
 AOI21xp33_ASAP7_75t_R n_1724 (.A1(n_1498_o_0),
    .A2(n_1511_o_0),
    .B(n_1661_o_0),
    .Y(n_1724_o_0));
 NAND3xp33_ASAP7_75t_R n_1725 (.A(n_1518_o_0),
    .B(n_1537_o_0),
    .C(n_1475_o_0),
    .Y(n_1725_o_0));
 OAI31xp33_ASAP7_75t_R n_1726 (.A1(n_1449_o_0),
    .A2(n_1725_o_0),
    .A3(n_1426_o_0),
    .B(n_1484_o_0),
    .Y(n_1726_o_0));
 AO21x1_ASAP7_75t_R n_1727 (.A1(n_1723_o_0),
    .A2(n_1724_o_0),
    .B(n_1726_o_0),
    .Y(n_1727_o_0));
 OAI211xp5_ASAP7_75t_R n_1728 (.A1(n_1406_o_0),
    .A2(n_1414_o_0),
    .B(n_1562_o_0),
    .C(n_1449_o_0),
    .Y(n_1728_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1729 (.A1(n_1527_o_0),
    .A2(n_1529_o_0),
    .B(n_1449_o_0),
    .C(n_1728_o_0),
    .Y(n_1729_o_0));
 NOR3xp33_ASAP7_75t_R n_1730 (.A(n_1729_o_0),
    .B(n_1496_o_0),
    .C(n_1400_o_0),
    .Y(n_1730_o_0));
 OAI21xp33_ASAP7_75t_R n_1731 (.A1(n_1727_o_0),
    .A2(n_1730_o_0),
    .B(n_1347_o_0),
    .Y(n_1731_o_0));
 AOI21xp33_ASAP7_75t_R n_1732 (.A1(n_1355_o_0),
    .A2(n_1722_o_0),
    .B(n_1731_o_0),
    .Y(n_1732_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_1733 (.A1(n_1695_o_0),
    .A2(n_1697_o_0),
    .B(n_1702_o_0),
    .C(n_1714_o_0),
    .D(n_1732_o_0),
    .Y(n_1733_o_0));
 OAI21xp33_ASAP7_75t_R n_1734 (.A1(n_1438_o_0),
    .A2(n_1561_o_0),
    .B(n_1629_o_0),
    .Y(n_1734_o_0));
 AOI21xp33_ASAP7_75t_R n_1735 (.A1(n_1496_o_0),
    .A2(n_1734_o_0),
    .B(n_1363_o_0),
    .Y(n_1735_o_0));
 INVx1_ASAP7_75t_R n_1736 (.A(n_1527_o_0),
    .Y(n_1736_o_0));
 AOI22xp33_ASAP7_75t_R n_1737 (.A1(n_1736_o_0),
    .A2(n_1466_o_0),
    .B1(net71),
    .B2(n_1467_o_0),
    .Y(n_1737_o_0));
 AOI21xp33_ASAP7_75t_R n_1738 (.A1(n_1496_o_0),
    .A2(n_1737_o_0),
    .B(n_1449_o_0),
    .Y(n_1738_o_0));
 AOI21xp33_ASAP7_75t_R n_1739 (.A1(n_1409_o_0),
    .A2(n_1415_o_0),
    .B(n_1542_o_0),
    .Y(n_1739_o_0));
 AOI21xp33_ASAP7_75t_R n_1740 (.A1(n_1508_o_0),
    .A2(n_1477_o_0),
    .B(n_1449_o_0),
    .Y(n_1740_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_1741 (.A1(net70),
    .A2(n_1387_o_0),
    .B(n_1404_o_0),
    .C(n_1518_o_0),
    .D(n_1363_o_0),
    .Y(n_1741_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1742 (.A1(net20),
    .A2(n_1739_o_0),
    .B(n_1740_o_0),
    .C(n_1741_o_0),
    .Y(n_1742_o_0));
 NAND2xp33_ASAP7_75t_R n_1743 (.A(n_1426_o_0),
    .B(n_1742_o_0),
    .Y(n_1743_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1744 (.A1(n_1735_o_0),
    .A2(n_1738_o_0),
    .B(n_1743_o_0),
    .C(n_1484_o_0),
    .Y(n_1744_o_0));
 AOI21xp33_ASAP7_75t_R n_1745 (.A1(n_1511_o_0),
    .A2(n_1435_o_0),
    .B(n_1363_o_0),
    .Y(n_1745_o_0));
 NAND3xp33_ASAP7_75t_R n_1746 (.A(n_1461_o_0),
    .B(n_1447_o_0),
    .C(net70),
    .Y(n_1746_o_0));
 OAI311xp33_ASAP7_75t_R n_1747 (.A1(n_1501_o_0),
    .A2(n_1669_o_0),
    .A3(net20),
    .B1(n_1363_o_0),
    .C1(n_1746_o_0),
    .Y(n_1747_o_0));
 INVx1_ASAP7_75t_R n_1748 (.A(n_1747_o_0),
    .Y(n_1748_o_0));
 AOI31xp33_ASAP7_75t_R n_1749 (.A1(n_1437_o_0),
    .A2(n_1518_o_0),
    .A3(n_1745_o_0),
    .B(n_1748_o_0),
    .Y(n_1749_o_0));
 INVx1_ASAP7_75t_R n_1750 (.A(n_1645_o_0),
    .Y(n_1750_o_0));
 NAND2xp33_ASAP7_75t_R n_1751 (.A(n_1363_o_0),
    .B(n_1566_o_0),
    .Y(n_1751_o_0));
 OAI32xp33_ASAP7_75t_R n_1752 (.A1(n_1489_o_0),
    .A2(n_1750_o_0),
    .A3(n_1363_o_0),
    .B1(n_1751_o_0),
    .B2(n_1562_o_0),
    .Y(n_1752_o_0));
 AOI21xp33_ASAP7_75t_R n_1753 (.A1(n_1484_o_0),
    .A2(n_1752_o_0),
    .B(n_1426_o_0),
    .Y(n_1753_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1754 (.A1(n_1355_o_0),
    .A2(n_1749_o_0),
    .B(n_1426_o_0),
    .C(n_1753_o_0),
    .Y(n_1754_o_0));
 AO21x1_ASAP7_75t_R n_1755 (.A1(n_1626_o_0),
    .A2(n_1581_o_0),
    .B(n_1496_o_0),
    .Y(n_1755_o_0));
 INVx1_ASAP7_75t_R n_1756 (.A(n_1478_o_0),
    .Y(n_1756_o_0));
 OAI21xp33_ASAP7_75t_R n_1757 (.A1(n_1410_o_0),
    .A2(n_1414_o_0),
    .B(n_1408_o_0),
    .Y(n_1757_o_0));
 OAI21xp33_ASAP7_75t_R n_1758 (.A1(n_1756_o_0),
    .A2(n_1644_o_0),
    .B(n_1757_o_0),
    .Y(n_1758_o_0));
 AOI21xp33_ASAP7_75t_R n_1759 (.A1(n_1496_o_0),
    .A2(n_1758_o_0),
    .B(n_1449_o_0),
    .Y(n_1759_o_0));
 OAI21xp33_ASAP7_75t_R n_1760 (.A1(net28),
    .A2(n_1388_o_0),
    .B(n_1407_o_0),
    .Y(n_1760_o_0));
 OAI21xp33_ASAP7_75t_R n_1761 (.A1(n_1760_o_0),
    .A2(n_1418_o_0),
    .B(n_1429_o_0),
    .Y(n_1761_o_0));
 OAI211xp5_ASAP7_75t_R n_1762 (.A1(n_1409_o_0),
    .A2(net20),
    .B(n_1723_o_0),
    .C(n_1760_o_0),
    .Y(n_1762_o_0));
 OAI21xp33_ASAP7_75t_R n_1763 (.A1(n_1560_o_0),
    .A2(n_1761_o_0),
    .B(n_1762_o_0),
    .Y(n_1763_o_0));
 AOI21xp33_ASAP7_75t_R n_1764 (.A1(n_1755_o_0),
    .A2(n_1759_o_0),
    .B(n_1763_o_0),
    .Y(n_1764_o_0));
 OAI21xp33_ASAP7_75t_R n_1765 (.A1(n_1760_o_0),
    .A2(n_1644_o_0),
    .B(n_1496_o_0),
    .Y(n_1765_o_0));
 AOI21xp33_ASAP7_75t_R n_1766 (.A1(n_1430_o_0),
    .A2(n_1447_o_0),
    .B(n_1496_o_0),
    .Y(n_1766_o_0));
 OAI21xp33_ASAP7_75t_R n_1767 (.A1(n_1561_o_0),
    .A2(n_1418_o_0),
    .B(n_1766_o_0),
    .Y(n_1767_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1768 (.A1(n_1410_o_0),
    .A2(n_1661_o_0),
    .B(n_1765_o_0),
    .C(n_1767_o_0),
    .Y(n_1768_o_0));
 OAI21xp33_ASAP7_75t_R n_1769 (.A1(n_1510_o_0),
    .A2(n_1669_o_0),
    .B(n_1399_o_0),
    .Y(n_1769_o_0));
 OAI22xp33_ASAP7_75t_R n_1770 (.A1(n_1497_o_0),
    .A2(n_1499_o_0),
    .B1(net13),
    .B2(n_1389_o_0),
    .Y(n_1770_o_0));
 NOR2xp33_ASAP7_75t_R n_1771 (.A(n_1363_o_0),
    .B(n_1496_o_0),
    .Y(n_1771_o_0));
 AOI22xp33_ASAP7_75t_R n_1772 (.A1(n_1769_o_0),
    .A2(n_1723_o_0),
    .B1(n_1770_o_0),
    .B2(n_1771_o_0),
    .Y(n_1772_o_0));
 OAI211xp5_ASAP7_75t_R n_1773 (.A1(n_1768_o_0),
    .A2(n_1449_o_0),
    .B(n_1484_o_0),
    .C(n_1772_o_0),
    .Y(n_1773_o_0));
 OAI211xp5_ASAP7_75t_R n_1774 (.A1(n_1764_o_0),
    .A2(n_1484_o_0),
    .B(n_1347_o_0),
    .C(n_1773_o_0),
    .Y(n_1774_o_0));
 OAI31xp33_ASAP7_75t_R n_1775 (.A1(n_1744_o_0),
    .A2(n_1754_o_0),
    .A3(n_1347_o_0),
    .B(n_1774_o_0),
    .Y(n_1775_o_0));
 AOI21xp33_ASAP7_75t_R n_1776 (.A1(n_1417_o_0),
    .A2(n_1489_o_0),
    .B(n_1449_o_0),
    .Y(n_1776_o_0));
 OAI21xp33_ASAP7_75t_R n_1777 (.A1(net13),
    .A2(n_1567_o_0),
    .B(n_1776_o_0),
    .Y(n_1777_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1778 (.A1(n_1436_o_0),
    .A2(n_1414_o_0),
    .B(n_1478_o_0),
    .C(n_1363_o_0),
    .Y(n_1778_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1779 (.A1(n_1404_o_0),
    .A2(net99),
    .B(n_1545_o_0),
    .C(n_1778_o_0),
    .Y(n_1779_o_0));
 AOI311xp33_ASAP7_75t_R n_1780 (.A1(n_1463_o_0),
    .A2(n_1461_o_0),
    .A3(net71),
    .B(n_1363_o_0),
    .C(n_1426_o_0),
    .Y(n_1780_o_0));
 OAI21xp33_ASAP7_75t_R n_1781 (.A1(n_1372_o_0),
    .A2(n_1409_o_0),
    .B(n_1446_o_0),
    .Y(n_1781_o_0));
 AOI211xp5_ASAP7_75t_R n_1782 (.A1(n_1781_o_0),
    .A2(n_1709_o_0),
    .B(n_1449_o_0),
    .C(n_1426_o_0),
    .Y(n_1782_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_1783 (.A1(n_1528_o_0),
    .A2(n_1415_o_0),
    .B(n_1497_o_0),
    .C(n_1780_o_0),
    .D(n_1782_o_0),
    .Y(n_1783_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1784 (.A1(n_1777_o_0),
    .A2(n_1779_o_0),
    .B(n_1496_o_0),
    .C(n_1783_o_0),
    .Y(n_1784_o_0));
 AOI21xp33_ASAP7_75t_R n_1785 (.A1(n_1723_o_0),
    .A2(n_1615_o_0),
    .B(n_1521_o_0),
    .Y(n_1785_o_0));
 NAND4xp25_ASAP7_75t_R n_1786 (.A(n_1717_o_0),
    .B(n_1541_o_0),
    .C(n_1496_o_0),
    .D(n_1363_o_0),
    .Y(n_1786_o_0));
 OAI211xp5_ASAP7_75t_R n_1787 (.A1(n_1581_o_0),
    .A2(n_1528_o_0),
    .B(n_1532_o_0),
    .C(n_1363_o_0),
    .Y(n_1787_o_0));
 NAND2xp33_ASAP7_75t_R n_1788 (.A(n_1380_o_0),
    .B(net28),
    .Y(n_1788_o_0));
 AOI211xp5_ASAP7_75t_R n_1789 (.A1(n_1430_o_0),
    .A2(n_1447_o_0),
    .B(n_1496_o_0),
    .C(n_1363_o_0),
    .Y(n_1789_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1790 (.A1(n_1788_o_0),
    .A2(n_1555_o_0),
    .B(net20),
    .C(n_1789_o_0),
    .Y(n_1790_o_0));
 NAND4xp25_ASAP7_75t_R n_1791 (.A(n_1785_o_0),
    .B(n_1786_o_0),
    .C(n_1787_o_0),
    .D(n_1790_o_0),
    .Y(n_1791_o_0));
 OAI21xp33_ASAP7_75t_R n_1792 (.A1(n_1347_o_0),
    .A2(n_1784_o_0),
    .B(n_1791_o_0),
    .Y(n_1792_o_0));
 NOR2xp33_ASAP7_75t_R n_1793 (.A(n_1484_o_0),
    .B(n_1792_o_0),
    .Y(n_1793_o_0));
 OAI21xp33_ASAP7_75t_R n_1794 (.A1(n_1510_o_0),
    .A2(n_1418_o_0),
    .B(n_1496_o_0),
    .Y(n_1794_o_0));
 AOI21xp33_ASAP7_75t_R n_1795 (.A1(n_1500_o_0),
    .A2(net71),
    .B(n_1705_o_0),
    .Y(n_1795_o_0));
 OAI21xp33_ASAP7_75t_R n_1796 (.A1(n_1464_o_0),
    .A2(n_1795_o_0),
    .B(n_1426_o_0),
    .Y(n_1796_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1797 (.A1(n_1556_o_0),
    .A2(net71),
    .B(n_1794_o_0),
    .C(n_1796_o_0),
    .Y(n_1797_o_0));
 OA21x2_ASAP7_75t_R n_1798 (.A1(n_1416_o_0),
    .A2(n_1414_o_0),
    .B(n_1430_o_0),
    .Y(n_1798_o_0));
 AOI31xp33_ASAP7_75t_R n_1799 (.A1(n_1463_o_0),
    .A2(n_1500_o_0),
    .A3(net71),
    .B(n_1798_o_0),
    .Y(n_1799_o_0));
 AOI211xp5_ASAP7_75t_R n_1800 (.A1(n_1409_o_0),
    .A2(net99),
    .B(net44),
    .C(n_1507_o_0),
    .Y(n_1800_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1801 (.A1(n_1478_o_0),
    .A2(n_1800_o_0),
    .B(n_1496_o_0),
    .C(n_1363_o_0),
    .Y(n_1801_o_0));
 OAI21xp33_ASAP7_75t_R n_1802 (.A1(n_1496_o_0),
    .A2(n_1799_o_0),
    .B(n_1801_o_0),
    .Y(n_1802_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1803 (.A1(n_1449_o_0),
    .A2(n_1797_o_0),
    .B(n_1802_o_0),
    .C(n_1521_o_0),
    .Y(n_1803_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1804 (.A1(n_1436_o_0),
    .A2(n_1452_o_0),
    .B(n_1705_o_0),
    .C(n_1447_o_0),
    .Y(n_1804_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1805 (.A1(n_1380_o_0),
    .A2(n_1387_o_0),
    .B(n_1656_o_0),
    .C(n_1804_o_0),
    .Y(n_1805_o_0));
 OAI211xp5_ASAP7_75t_R n_1806 (.A1(n_1467_o_0),
    .A2(n_1497_o_0),
    .B(n_1645_o_0),
    .C(n_1363_o_0),
    .Y(n_1806_o_0));
 OAI211xp5_ASAP7_75t_R n_1807 (.A1(n_1805_o_0),
    .A2(n_1363_o_0),
    .B(n_1496_o_0),
    .C(n_1806_o_0),
    .Y(n_1807_o_0));
 AOI21xp33_ASAP7_75t_R n_1808 (.A1(n_1555_o_0),
    .A2(n_1477_o_0),
    .B(net44),
    .Y(n_1808_o_0));
 OAI21xp33_ASAP7_75t_R n_1809 (.A1(n_1380_o_0),
    .A2(net71),
    .B(n_1449_o_0),
    .Y(n_1809_o_0));
 NAND2xp33_ASAP7_75t_R n_1810 (.A(n_1436_o_0),
    .B(n_1661_o_0),
    .Y(n_1810_o_0));
 NAND4xp25_ASAP7_75t_R n_1811 (.A(n_1649_o_0),
    .B(n_1810_o_0),
    .C(n_1475_o_0),
    .D(n_1363_o_0),
    .Y(n_1811_o_0));
 OAI211xp5_ASAP7_75t_R n_1812 (.A1(n_1808_o_0),
    .A2(n_1809_o_0),
    .B(n_1811_o_0),
    .C(n_1426_o_0),
    .Y(n_1812_o_0));
 AOI21xp33_ASAP7_75t_R n_1813 (.A1(n_1807_o_0),
    .A2(n_1812_o_0),
    .B(n_1347_o_0),
    .Y(n_1813_o_0));
 OAI211xp5_ASAP7_75t_R n_1814 (.A1(n_1784_o_0),
    .A2(n_1347_o_0),
    .B(n_1355_o_0),
    .C(n_1791_o_0),
    .Y(n_1814_o_0));
 OAI211xp5_ASAP7_75t_R n_1815 (.A1(n_1803_o_0),
    .A2(n_1813_o_0),
    .B(n_1814_o_0),
    .C(n_1484_o_0),
    .Y(n_1815_o_0));
 OAI21xp33_ASAP7_75t_R n_1816 (.A1(n_1484_o_0),
    .A2(n_1793_o_0),
    .B(n_1815_o_0),
    .Y(n_1816_o_0));
 INVx1_ASAP7_75t_R n_1817 (.A(n_1475_o_0),
    .Y(n_1817_o_0));
 AOI21xp33_ASAP7_75t_R n_1818 (.A1(n_1675_o_0),
    .A2(net71),
    .B(n_1817_o_0),
    .Y(n_1818_o_0));
 NAND3xp33_ASAP7_75t_R n_1819 (.A(n_1388_o_0),
    .B(net20),
    .C(net28),
    .Y(n_1819_o_0));
 OAI31xp33_ASAP7_75t_R n_1820 (.A1(net71),
    .A2(n_1487_o_0),
    .A3(n_1567_o_0),
    .B(n_1363_o_0),
    .Y(n_1820_o_0));
 AOI21xp33_ASAP7_75t_R n_1821 (.A1(n_1628_o_0),
    .A2(n_1447_o_0),
    .B(n_1820_o_0),
    .Y(n_1821_o_0));
 AOI311xp33_ASAP7_75t_R n_1822 (.A1(n_1449_o_0),
    .A2(n_1818_o_0),
    .A3(n_1819_o_0),
    .B(n_1496_o_0),
    .C(n_1821_o_0),
    .Y(n_1822_o_0));
 AOI21xp33_ASAP7_75t_R n_1823 (.A1(net20),
    .A2(n_1416_o_0),
    .B(n_1808_o_0),
    .Y(n_1823_o_0));
 AOI211xp5_ASAP7_75t_R n_1824 (.A1(net70),
    .A2(n_1387_o_0),
    .B(net99),
    .C(n_1380_o_0),
    .Y(n_1824_o_0));
 NOR3xp33_ASAP7_75t_R n_1825 (.A(n_1574_o_0),
    .B(n_1824_o_0),
    .C(n_1363_o_0),
    .Y(n_1825_o_0));
 AOI211xp5_ASAP7_75t_R n_1826 (.A1(n_1363_o_0),
    .A2(n_1823_o_0),
    .B(n_1825_o_0),
    .C(n_1426_o_0),
    .Y(n_1826_o_0));
 NOR3xp33_ASAP7_75t_R n_1827 (.A(n_1822_o_0),
    .B(n_1355_o_0),
    .C(n_1826_o_0),
    .Y(n_1827_o_0));
 OAI21xp33_ASAP7_75t_R n_1828 (.A1(n_1406_o_0),
    .A2(n_1414_o_0),
    .B(n_1408_o_0),
    .Y(n_1828_o_0));
 OAI31xp33_ASAP7_75t_R n_1829 (.A1(net71),
    .A2(n_1464_o_0),
    .A3(n_1567_o_0),
    .B(n_1828_o_0),
    .Y(n_1829_o_0));
 NAND3xp33_ASAP7_75t_R n_1830 (.A(n_1455_o_0),
    .B(n_1518_o_0),
    .C(n_1537_o_0),
    .Y(n_1830_o_0));
 AOI21xp33_ASAP7_75t_R n_1831 (.A1(n_1426_o_0),
    .A2(n_1830_o_0),
    .B(n_1449_o_0),
    .Y(n_1831_o_0));
 OAI21xp33_ASAP7_75t_R n_1832 (.A1(n_1829_o_0),
    .A2(n_1426_o_0),
    .B(n_1831_o_0),
    .Y(n_1832_o_0));
 NAND2xp33_ASAP7_75t_R n_1833 (.A(net44),
    .B(n_1431_o_0),
    .Y(n_1833_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1834 (.A1(n_1539_o_0),
    .A2(net20),
    .B(n_1833_o_0),
    .C(n_1412_o_0),
    .Y(n_1834_o_0));
 OAI31xp33_ASAP7_75t_R n_1835 (.A1(net99),
    .A2(n_1473_o_0),
    .A3(net71),
    .B(n_1771_o_0),
    .Y(n_1835_o_0));
 AOI21xp33_ASAP7_75t_R n_1836 (.A1(net71),
    .A2(n_1388_o_0),
    .B(n_1835_o_0),
    .Y(n_1836_o_0));
 AOI21xp33_ASAP7_75t_R n_1837 (.A1(n_1723_o_0),
    .A2(n_1834_o_0),
    .B(n_1836_o_0),
    .Y(n_1837_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1838 (.A1(n_1832_o_0),
    .A2(n_1837_o_0),
    .B(n_1484_o_0),
    .C(n_1521_o_0),
    .Y(n_1838_o_0));
 OAI21xp33_ASAP7_75t_R n_1839 (.A1(net13),
    .A2(n_1462_o_0),
    .B(n_1363_o_0),
    .Y(n_1839_o_0));
 AOI21xp33_ASAP7_75t_R n_1840 (.A1(n_1488_o_0),
    .A2(n_1478_o_0),
    .B(n_1839_o_0),
    .Y(n_1840_o_0));
 NOR2xp33_ASAP7_75t_R n_1841 (.A(net28),
    .B(net13),
    .Y(n_1841_o_0));
 AOI211xp5_ASAP7_75t_R n_1842 (.A1(n_1388_o_0),
    .A2(n_1841_o_0),
    .B(n_1655_o_0),
    .C(n_1363_o_0),
    .Y(n_1842_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1843 (.A1(n_1488_o_0),
    .A2(n_1430_o_0),
    .B(n_1600_o_0),
    .C(n_1771_o_0),
    .Y(n_1843_o_0));
 OAI31xp33_ASAP7_75t_R n_1844 (.A1(n_1426_o_0),
    .A2(n_1840_o_0),
    .A3(n_1842_o_0),
    .B(n_1843_o_0),
    .Y(n_1844_o_0));
 AOI22xp33_ASAP7_75t_R n_1845 (.A1(n_1628_o_0),
    .A2(n_1540_o_0),
    .B1(net20),
    .B2(n_1387_o_0),
    .Y(n_1845_o_0));
 NOR3xp33_ASAP7_75t_R n_1846 (.A(n_1845_o_0),
    .B(n_1449_o_0),
    .C(n_1496_o_0),
    .Y(n_1846_o_0));
 OAI22xp33_ASAP7_75t_R n_1847 (.A1(n_1643_o_0),
    .A2(n_1507_o_0),
    .B1(n_1553_o_0),
    .B2(net70),
    .Y(n_1847_o_0));
 AOI21xp33_ASAP7_75t_R n_1848 (.A1(net71),
    .A2(n_1687_o_0),
    .B(n_1363_o_0),
    .Y(n_1848_o_0));
 OAI31xp33_ASAP7_75t_R n_1849 (.A1(net71),
    .A2(n_1448_o_0),
    .A3(n_1515_o_0),
    .B(n_1848_o_0),
    .Y(n_1849_o_0));
 OAI211xp5_ASAP7_75t_R n_1850 (.A1(n_1847_o_0),
    .A2(n_1449_o_0),
    .B(n_1496_o_0),
    .C(n_1849_o_0),
    .Y(n_1850_o_0));
 NAND2xp33_ASAP7_75t_R n_1851 (.A(n_1388_o_0),
    .B(n_1661_o_0),
    .Y(n_1851_o_0));
 OAI31xp33_ASAP7_75t_R n_1852 (.A1(net71),
    .A2(n_1462_o_0),
    .A3(n_1507_o_0),
    .B(n_1851_o_0),
    .Y(n_1852_o_0));
 OAI211xp5_ASAP7_75t_R n_1853 (.A1(net71),
    .A2(n_1515_o_0),
    .B(n_1717_o_0),
    .C(n_1449_o_0),
    .Y(n_1853_o_0));
 OAI311xp33_ASAP7_75t_R n_1854 (.A1(n_1458_o_0),
    .A2(n_1852_o_0),
    .A3(n_1449_o_0),
    .B1(n_1853_o_0),
    .C1(n_1426_o_0),
    .Y(n_1854_o_0));
 NAND3xp33_ASAP7_75t_R n_1855 (.A(n_1850_o_0),
    .B(n_1854_o_0),
    .C(n_1484_o_0),
    .Y(n_1855_o_0));
 OAI311xp33_ASAP7_75t_R n_1856 (.A1(n_1844_o_0),
    .A2(n_1846_o_0),
    .A3(n_1484_o_0),
    .B1(n_1347_o_0),
    .C1(n_1855_o_0),
    .Y(n_1856_o_0));
 OAI21xp33_ASAP7_75t_R n_1857 (.A1(n_1827_o_0),
    .A2(n_1838_o_0),
    .B(n_1856_o_0),
    .Y(n_1857_o_0));
 INVx1_ASAP7_75t_R n_1858 (.A(_00963_),
    .Y(n_1858_o_0));
 XNOR2xp5_ASAP7_75t_R n_1859 (.A(_00431_),
    .B(_00867_),
    .Y(n_1859_o_0));
 XNOR2xp5_ASAP7_75t_R n_1860 (.A(_00899_),
    .B(n_1859_o_0),
    .Y(n_1860_o_0));
 INVx1_ASAP7_75t_R n_1861 (.A(n_1860_o_0),
    .Y(n_1861_o_0));
 XNOR2xp5_ASAP7_75t_R n_1862 (.A(_00931_),
    .B(n_1861_o_0),
    .Y(n_1862_o_0));
 NOR2xp33_ASAP7_75t_R n_1863 (.A(n_1858_o_0),
    .B(n_1862_o_0),
    .Y(n_1863_o_0));
 AOI211xp5_ASAP7_75t_R n_1864 (.A1(n_1858_o_0),
    .A2(n_1862_o_0),
    .B(n_1863_o_0),
    .C(ld),
    .Y(n_1864_o_0));
 AOI21xp33_ASAP7_75t_R n_1865 (.A1(key[7]),
    .A2(ld),
    .B(n_1864_o_0),
    .Y(n_1865_o_0));
 XNOR2xp5_ASAP7_75t_R n_1866 (.A(_00430_),
    .B(_00866_),
    .Y(n_1866_o_0));
 XNOR2xp5_ASAP7_75t_R n_1867 (.A(_00898_),
    .B(n_1866_o_0),
    .Y(n_1867_o_0));
 INVx1_ASAP7_75t_R n_1868 (.A(n_1867_o_0),
    .Y(n_1868_o_0));
 XNOR2xp5_ASAP7_75t_R n_1869 (.A(_00930_),
    .B(n_1868_o_0),
    .Y(n_1869_o_0));
 XNOR2xp5_ASAP7_75t_R n_1870 (.A(_00962_),
    .B(n_1869_o_0),
    .Y(n_1870_o_0));
 OR2x2_ASAP7_75t_R n_1871 (.A(key[6]),
    .B(n_827_o_0),
    .Y(n_1871_o_0));
 OAI21xp33_ASAP7_75t_R n_1872 (.A1(ld),
    .A2(n_1870_o_0),
    .B(n_1871_o_0),
    .Y(n_1872_o_0));
 INVx1_ASAP7_75t_R n_1873 (.A(n_1872_o_0),
    .Y(n_1873_o_0));
 XOR2xp5_ASAP7_75t_R n_1874 (.A(_00429_),
    .B(_00865_),
    .Y(n_1874_o_0));
 XNOR2xp5_ASAP7_75t_R n_1875 (.A(_00897_),
    .B(n_1874_o_0),
    .Y(n_1875_o_0));
 XNOR2xp5_ASAP7_75t_R n_1876 (.A(_00929_),
    .B(n_1875_o_0),
    .Y(n_1876_o_0));
 INVx1_ASAP7_75t_R n_1877 (.A(_00961_),
    .Y(n_1877_o_0));
 NOR2xp33_ASAP7_75t_R n_1878 (.A(n_1877_o_0),
    .B(n_1876_o_0),
    .Y(n_1878_o_0));
 NOR2xp33_ASAP7_75t_R n_1879 (.A(key[5]),
    .B(n_827_o_0),
    .Y(n_1879_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_1880 (.A1(n_1876_o_0),
    .A2(n_1877_o_0),
    .B(n_1878_o_0),
    .C(n_827_o_0),
    .D(n_1879_o_0),
    .Y(n_1880_o_0));
 XOR2xp5_ASAP7_75t_R n_1881 (.A(_00428_),
    .B(_00864_),
    .Y(n_1881_o_0));
 XNOR2xp5_ASAP7_75t_R n_1882 (.A(_00896_),
    .B(n_1881_o_0),
    .Y(n_1882_o_0));
 INVx1_ASAP7_75t_R n_1883 (.A(_00928_),
    .Y(n_1883_o_0));
 NAND2xp33_ASAP7_75t_R n_1884 (.A(n_1883_o_0),
    .B(n_1882_o_0),
    .Y(n_1884_o_0));
 OAI21xp33_ASAP7_75t_R n_1885 (.A1(n_1882_o_0),
    .A2(n_1883_o_0),
    .B(n_1884_o_0),
    .Y(n_1885_o_0));
 NAND2xp33_ASAP7_75t_R n_1886 (.A(_00960_),
    .B(n_1885_o_0),
    .Y(n_1886_o_0));
 INVx1_ASAP7_75t_R n_1887 (.A(_00960_),
    .Y(n_1887_o_0));
 OAI211xp5_ASAP7_75t_R n_1888 (.A1(n_1883_o_0),
    .A2(n_1882_o_0),
    .B(n_1884_o_0),
    .C(n_1887_o_0),
    .Y(n_1888_o_0));
 AND2x2_ASAP7_75t_R n_1889 (.A(key[4]),
    .B(ld),
    .Y(n_1889_o_0));
 AOI31xp67_ASAP7_75t_R n_1890 (.A1(n_827_o_0),
    .A2(n_1886_o_0),
    .A3(n_1888_o_0),
    .B(n_1889_o_0),
    .Y(n_1890_o_0));
 XNOR2xp5_ASAP7_75t_R n_1891 (.A(_00423_),
    .B(_00862_),
    .Y(n_1891_o_0));
 AND2x2_ASAP7_75t_R n_1892 (.A(n_827_o_0),
    .B(n_1891_o_0),
    .Y(n_1892_o_0));
 XOR2xp5_ASAP7_75t_R n_1893 (.A(_00926_),
    .B(_00958_),
    .Y(n_1893_o_0));
 XNOR2xp5_ASAP7_75t_R n_1894 (.A(_00894_),
    .B(n_1893_o_0),
    .Y(n_1894_o_0));
 NAND2xp33_ASAP7_75t_R n_1895 (.A(n_1892_o_0),
    .B(n_1894_o_0),
    .Y(n_1895_o_0));
 NOR3xp33_ASAP7_75t_R n_1896 (.A(n_1894_o_0),
    .B(n_1891_o_0),
    .C(ld),
    .Y(n_1896_o_0));
 AOI21xp33_ASAP7_75t_R n_1897 (.A1(key[2]),
    .A2(ld),
    .B(n_1896_o_0),
    .Y(n_1897_o_0));
 NAND2x1p5_ASAP7_75t_R n_1898 (.A(n_1895_o_0),
    .B(n_1897_o_0),
    .Y(n_1898_o_0));
 XNOR2xp5_ASAP7_75t_R n_1899 (.A(_00924_),
    .B(_00956_),
    .Y(n_1899_o_0));
 XNOR2xp5_ASAP7_75t_R n_1900 (.A(_00425_),
    .B(_00860_),
    .Y(n_1900_o_0));
 NAND2xp33_ASAP7_75t_R n_1901 (.A(_00892_),
    .B(n_1900_o_0),
    .Y(n_1901_o_0));
 OAI21xp33_ASAP7_75t_R n_1902 (.A1(_00892_),
    .A2(n_1900_o_0),
    .B(n_1901_o_0),
    .Y(n_1902_o_0));
 XNOR2xp5_ASAP7_75t_R n_1903 (.A(n_1899_o_0),
    .B(n_1902_o_0),
    .Y(n_1903_o_0));
 NOR2xp33_ASAP7_75t_R n_1904 (.A(_00925_),
    .B(_00957_),
    .Y(n_1904_o_0));
 XNOR2xp5_ASAP7_75t_R n_1905 (.A(_00426_),
    .B(_00861_),
    .Y(n_1905_o_0));
 NAND2xp33_ASAP7_75t_R n_1906 (.A(_00893_),
    .B(n_1905_o_0),
    .Y(n_1906_o_0));
 OAI21xp33_ASAP7_75t_R n_1907 (.A1(_00893_),
    .A2(n_1905_o_0),
    .B(n_1906_o_0),
    .Y(n_1907_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1908 (.A1(_00925_),
    .A2(_00957_),
    .B(n_1904_o_0),
    .C(n_1907_o_0),
    .Y(n_1908_o_0));
 AOI21xp33_ASAP7_75t_R n_1909 (.A1(_00925_),
    .A2(_00957_),
    .B(n_1904_o_0),
    .Y(n_1909_o_0));
 OAI211xp5_ASAP7_75t_R n_1910 (.A1(_00893_),
    .A2(n_1905_o_0),
    .B(n_1906_o_0),
    .C(n_1909_o_0),
    .Y(n_1910_o_0));
 AND2x2_ASAP7_75t_R n_1911 (.A(key[1]),
    .B(ld),
    .Y(n_1911_o_0));
 AOI31xp33_ASAP7_75t_R n_1912 (.A1(n_827_o_0),
    .A2(n_1908_o_0),
    .A3(n_1910_o_0),
    .B(n_1911_o_0),
    .Y(n_1912_o_0));
 NOR2xp33_ASAP7_75t_R n_1913 (.A(key[0]),
    .B(n_827_o_0),
    .Y(n_1913_o_0));
 AOI211xp5_ASAP7_75t_R n_1914 (.A1(n_1903_o_0),
    .A2(n_827_o_0),
    .B(n_1912_o_0),
    .C(n_1913_o_0),
    .Y(n_1914_o_0));
 INVx1_ASAP7_75t_R n_1915 (.A(n_1914_o_0),
    .Y(n_1915_o_0));
 AOI21x1_ASAP7_75t_R n_1916 (.A1(n_827_o_0),
    .A2(n_1903_o_0),
    .B(n_1913_o_0),
    .Y(n_1916_o_0));
 INVx1_ASAP7_75t_R n_1917 (.A(n_1916_o_0),
    .Y(n_1917_o_0));
 NOR2xp33_ASAP7_75t_R n_1918 (.A(n_1898_o_0),
    .B(n_1917_o_0),
    .Y(n_1918_o_0));
 XOR2xp5_ASAP7_75t_R n_1919 (.A(_00427_),
    .B(_00863_),
    .Y(n_1919_o_0));
 XNOR2xp5_ASAP7_75t_R n_1920 (.A(_00895_),
    .B(n_1919_o_0),
    .Y(n_1920_o_0));
 NOR2xp33_ASAP7_75t_R n_1921 (.A(_00927_),
    .B(n_1920_o_0),
    .Y(n_1921_o_0));
 INVx1_ASAP7_75t_R n_1922 (.A(_00959_),
    .Y(n_1922_o_0));
 AOI211xp5_ASAP7_75t_R n_1923 (.A1(_00927_),
    .A2(n_1920_o_0),
    .B(n_1921_o_0),
    .C(n_1922_o_0),
    .Y(n_1923_o_0));
 NAND2xp33_ASAP7_75t_R n_1924 (.A(_00927_),
    .B(n_1920_o_0),
    .Y(n_1924_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_1925 (.A1(_00927_),
    .A2(n_1920_o_0),
    .B(n_1924_o_0),
    .C(_00959_),
    .Y(n_1925_o_0));
 NAND2xp33_ASAP7_75t_R n_1926 (.A(key[3]),
    .B(ld),
    .Y(n_1926_o_0));
 OAI31xp67_ASAP7_75t_R n_1927 (.A1(n_1925_o_0),
    .A2(n_1923_o_0),
    .A3(ld),
    .B(n_1926_o_0),
    .Y(n_1927_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1928 (.A1(n_1898_o_0),
    .A2(n_1915_o_0),
    .B(n_1918_o_0),
    .C(n_1927_o_0),
    .Y(n_1928_o_0));
 INVx1_ASAP7_75t_R n_1929 (.A(n_1928_o_0),
    .Y(n_1929_o_0));
 INVx1_ASAP7_75t_R n_1930 (.A(n_1895_o_0),
    .Y(n_1930_o_0));
 AO21x1_ASAP7_75t_R n_1931 (.A1(key[2]),
    .A2(ld),
    .B(n_1896_o_0),
    .Y(n_1931_o_0));
 NOR2x1_ASAP7_75t_R n_1932 (.A(n_1930_o_0),
    .B(n_1931_o_0),
    .Y(n_1932_o_0));
 AOI211xp5_ASAP7_75t_R n_1933 (.A1(n_1903_o_0),
    .A2(n_827_o_0),
    .B(n_1912_o_0),
    .C(n_1913_o_0),
    .Y(n_1933_o_0));
 AOI21xp5_ASAP7_75t_R n_1934 (.A1(n_1912_o_0),
    .A2(n_1917_o_0),
    .B(n_1933_o_0),
    .Y(n_1934_o_0));
 OAI21xp33_ASAP7_75t_R n_1935 (.A1(n_1932_o_0),
    .A2(n_1934_o_0),
    .B(n_1927_o_0),
    .Y(n_1935_o_0));
 NAND2xp5_ASAP7_75t_R n_1936 (.A(n_1912_o_0),
    .B(n_1916_o_0),
    .Y(n_1936_o_0));
 INVx1_ASAP7_75t_R n_1937 (.A(n_1936_o_0),
    .Y(n_1937_o_0));
 INVx2_ASAP7_75t_R n_1938 (.A(n_1927_o_0),
    .Y(n_1938_o_0));
 NAND3xp33_ASAP7_75t_R n_1939 (.A(n_1937_o_0),
    .B(n_1898_o_0),
    .C(n_1938_o_0),
    .Y(n_1939_o_0));
 AOI21xp33_ASAP7_75t_R n_1940 (.A1(n_1935_o_0),
    .A2(n_1939_o_0),
    .B(n_1890_o_0),
    .Y(n_1940_o_0));
 AO31x2_ASAP7_75t_R n_1941 (.A1(n_1908_o_0),
    .A2(n_1910_o_0),
    .A3(n_827_o_0),
    .B(n_1911_o_0),
    .Y(n_1941_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1942 (.A1(n_1903_o_0),
    .A2(n_827_o_0),
    .B(n_1913_o_0),
    .C(n_1941_o_0),
    .Y(n_1942_o_0));
 NOR3xp33_ASAP7_75t_R n_1943 (.A(n_1927_o_0),
    .B(n_1898_o_0),
    .C(n_1942_o_0),
    .Y(n_1943_o_0));
 AOI211xp5_ASAP7_75t_R n_1944 (.A1(n_1890_o_0),
    .A2(n_1929_o_0),
    .B(n_1940_o_0),
    .C(n_1943_o_0),
    .Y(n_1944_o_0));
 NAND2xp33_ASAP7_75t_R n_1945 (.A(n_1898_o_0),
    .B(n_1917_o_0),
    .Y(n_1945_o_0));
 OAI211xp5_ASAP7_75t_R n_1946 (.A1(n_1898_o_0),
    .A2(n_1936_o_0),
    .B(n_1945_o_0),
    .C(net33),
    .Y(n_1946_o_0));
 INVx1_ASAP7_75t_R n_1947 (.A(n_1933_o_0),
    .Y(n_1947_o_0));
 OAI21xp33_ASAP7_75t_R n_1948 (.A1(n_1916_o_0),
    .A2(n_1941_o_0),
    .B(n_1947_o_0),
    .Y(n_1948_o_0));
 NAND2xp33_ASAP7_75t_R n_1949 (.A(n_1941_o_0),
    .B(n_1898_o_0),
    .Y(n_1949_o_0));
 OAI211xp5_ASAP7_75t_R n_1950 (.A1(n_1948_o_0),
    .A2(n_1898_o_0),
    .B(n_1938_o_0),
    .C(n_1949_o_0),
    .Y(n_1950_o_0));
 INVx1_ASAP7_75t_R n_1951 (.A(n_1890_o_0),
    .Y(n_1951_o_0));
 AOI21xp33_ASAP7_75t_R n_1952 (.A1(n_1946_o_0),
    .A2(n_1950_o_0),
    .B(n_1951_o_0),
    .Y(n_1952_o_0));
 INVx1_ASAP7_75t_R n_1953 (.A(n_1942_o_0),
    .Y(n_1953_o_0));
 OAI21xp33_ASAP7_75t_R n_1954 (.A1(n_1932_o_0),
    .A2(n_1953_o_0),
    .B(n_1927_o_0),
    .Y(n_1954_o_0));
 NOR2xp67_ASAP7_75t_R n_1955 (.A(n_1941_o_0),
    .B(n_1916_o_0),
    .Y(n_1955_o_0));
 NOR2xp33_ASAP7_75t_R n_1956 (.A(n_1898_o_0),
    .B(n_1955_o_0),
    .Y(n_1956_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1957 (.A1(n_1955_o_0),
    .A2(n_1898_o_0),
    .B(n_1956_o_0),
    .C(n_1938_o_0),
    .Y(n_1957_o_0));
 AOI21xp33_ASAP7_75t_R n_1958 (.A1(n_1954_o_0),
    .A2(n_1957_o_0),
    .B(n_1890_o_0),
    .Y(n_1958_o_0));
 OAI21xp33_ASAP7_75t_R n_1959 (.A1(n_1952_o_0),
    .A2(n_1958_o_0),
    .B(net31),
    .Y(n_1959_o_0));
 OAI21xp33_ASAP7_75t_R n_1960 (.A1(net31),
    .A2(n_1944_o_0),
    .B(n_1959_o_0),
    .Y(n_1960_o_0));
 OR2x2_ASAP7_75t_R n_1961 (.A(ld),
    .B(n_1870_o_0),
    .Y(n_1961_o_0));
 OAI21xp33_ASAP7_75t_R n_1962 (.A1(n_1930_o_0),
    .A2(n_1931_o_0),
    .B(n_1953_o_0),
    .Y(n_1962_o_0));
 OAI21xp33_ASAP7_75t_R n_1963 (.A1(n_1898_o_0),
    .A2(n_1936_o_0),
    .B(n_1938_o_0),
    .Y(n_1963_o_0));
 INVx1_ASAP7_75t_R n_1964 (.A(n_1963_o_0),
    .Y(n_1964_o_0));
 INVx1_ASAP7_75t_R n_1965 (.A(n_1955_o_0),
    .Y(n_1965_o_0));
 NOR3xp33_ASAP7_75t_R n_1966 (.A(n_1965_o_0),
    .B(n_1938_o_0),
    .C(n_1932_o_0),
    .Y(n_1966_o_0));
 AO21x1_ASAP7_75t_R n_1967 (.A1(n_1962_o_0),
    .A2(n_1964_o_0),
    .B(n_1966_o_0),
    .Y(n_1967_o_0));
 NAND2xp33_ASAP7_75t_R n_1968 (.A(n_1932_o_0),
    .B(n_1936_o_0),
    .Y(n_1968_o_0));
 NAND3xp33_ASAP7_75t_R n_1969 (.A(n_1968_o_0),
    .B(n_1962_o_0),
    .C(n_1927_o_0),
    .Y(n_1969_o_0));
 NAND3xp33_ASAP7_75t_R n_1970 (.A(n_1938_o_0),
    .B(n_1898_o_0),
    .C(n_1955_o_0),
    .Y(n_1970_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1971 (.A1(n_1969_o_0),
    .A2(n_1970_o_0),
    .B(n_1951_o_0),
    .C(n_1880_o_0),
    .Y(n_1971_o_0));
 AOI21xp33_ASAP7_75t_R n_1972 (.A1(net18),
    .A2(n_1967_o_0),
    .B(n_1971_o_0),
    .Y(n_1972_o_0));
 INVx1_ASAP7_75t_R n_1973 (.A(n_1949_o_0),
    .Y(n_1973_o_0));
 NOR2xp33_ASAP7_75t_R n_1974 (.A(n_1941_o_0),
    .B(n_1916_o_0),
    .Y(n_1974_o_0));
 OAI31xp33_ASAP7_75t_R n_1975 (.A1(n_1933_o_0),
    .A2(n_1974_o_0),
    .A3(n_1898_o_0),
    .B(n_1938_o_0),
    .Y(n_1975_o_0));
 OA21x2_ASAP7_75t_R n_1976 (.A1(n_1973_o_0),
    .A2(net4),
    .B(n_1975_o_0),
    .Y(n_1976_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_1977 (.A1(n_1965_o_0),
    .A2(n_1898_o_0),
    .B(n_1918_o_0),
    .C(n_1927_o_0),
    .Y(n_1977_o_0));
 NAND2xp33_ASAP7_75t_R n_1978 (.A(n_1916_o_0),
    .B(n_1932_o_0),
    .Y(n_1978_o_0));
 NAND3xp33_ASAP7_75t_R n_1979 (.A(n_1978_o_0),
    .B(n_1962_o_0),
    .C(net4),
    .Y(n_1979_o_0));
 AOI21xp33_ASAP7_75t_R n_1980 (.A1(n_1977_o_0),
    .A2(n_1979_o_0),
    .B(n_1951_o_0),
    .Y(n_1980_o_0));
 AOI211xp5_ASAP7_75t_R n_1981 (.A1(net17),
    .A2(n_1976_o_0),
    .B(n_1980_o_0),
    .C(n_1880_o_0),
    .Y(n_1981_o_0));
 AOI211xp5_ASAP7_75t_R n_1982 (.A1(n_1961_o_0),
    .A2(n_1871_o_0),
    .B(n_1972_o_0),
    .C(n_1981_o_0),
    .Y(n_1982_o_0));
 AOI21xp33_ASAP7_75t_R n_1983 (.A1(n_1873_o_0),
    .A2(n_1960_o_0),
    .B(n_1982_o_0),
    .Y(n_1983_o_0));
 NAND2xp33_ASAP7_75t_R n_1984 (.A(n_1932_o_0),
    .B(n_1953_o_0),
    .Y(n_1984_o_0));
 INVx1_ASAP7_75t_R n_1985 (.A(n_1954_o_0),
    .Y(n_1985_o_0));
 NOR2xp33_ASAP7_75t_R n_1986 (.A(n_1916_o_0),
    .B(n_1898_o_0),
    .Y(n_1986_o_0));
 OAI21xp33_ASAP7_75t_R n_1987 (.A1(net33),
    .A2(n_1986_o_0),
    .B(n_1890_o_0),
    .Y(n_1987_o_0));
 AOI21xp33_ASAP7_75t_R n_1988 (.A1(n_1984_o_0),
    .A2(n_1985_o_0),
    .B(n_1987_o_0),
    .Y(n_1988_o_0));
 NOR2xp33_ASAP7_75t_R n_1989 (.A(n_1914_o_0),
    .B(n_1898_o_0),
    .Y(n_1989_o_0));
 OAI21xp33_ASAP7_75t_R n_1990 (.A1(n_1932_o_0),
    .A2(n_1934_o_0),
    .B(n_1927_o_0),
    .Y(n_1990_o_0));
 OAI21xp33_ASAP7_75t_R n_1991 (.A1(n_1989_o_0),
    .A2(n_1990_o_0),
    .B(n_1951_o_0),
    .Y(n_1991_o_0));
 AOI31xp33_ASAP7_75t_R n_1992 (.A1(net8),
    .A2(n_1945_o_0),
    .A3(n_1984_o_0),
    .B(n_1991_o_0),
    .Y(n_1992_o_0));
 INVx2_ASAP7_75t_R n_1993 (.A(n_1880_o_0),
    .Y(n_1993_o_0));
 NOR2xp33_ASAP7_75t_R n_1994 (.A(n_1941_o_0),
    .B(n_1898_o_0),
    .Y(n_1994_o_0));
 INVx1_ASAP7_75t_R n_1995 (.A(n_1994_o_0),
    .Y(n_1995_o_0));
 OAI211xp5_ASAP7_75t_R n_1996 (.A1(n_1995_o_0),
    .A2(net33),
    .B(n_1928_o_0),
    .C(n_1970_o_0),
    .Y(n_1996_o_0));
 OAI211xp5_ASAP7_75t_R n_1997 (.A1(n_1932_o_0),
    .A2(n_1941_o_0),
    .B(net33),
    .C(n_1916_o_0),
    .Y(n_1997_o_0));
 NAND2xp33_ASAP7_75t_R n_1998 (.A(n_1912_o_0),
    .B(n_1898_o_0),
    .Y(n_1998_o_0));
 AOI31xp33_ASAP7_75t_R n_1999 (.A1(net4),
    .A2(n_1984_o_0),
    .A3(n_1998_o_0),
    .B(n_1890_o_0),
    .Y(n_1999_o_0));
 AOI21xp33_ASAP7_75t_R n_2000 (.A1(n_1997_o_0),
    .A2(n_1999_o_0),
    .B(net31),
    .Y(n_2000_o_0));
 OAI21xp33_ASAP7_75t_R n_2001 (.A1(net18),
    .A2(n_1996_o_0),
    .B(n_2000_o_0),
    .Y(n_2001_o_0));
 OAI31xp33_ASAP7_75t_R n_2002 (.A1(n_1988_o_0),
    .A2(n_1992_o_0),
    .A3(n_1993_o_0),
    .B(n_2001_o_0),
    .Y(n_2002_o_0));
 AOI21xp33_ASAP7_75t_R n_2003 (.A1(n_1898_o_0),
    .A2(n_1948_o_0),
    .B(n_1927_o_0),
    .Y(n_2003_o_0));
 OAI21xp33_ASAP7_75t_R n_2004 (.A1(n_1898_o_0),
    .A2(n_1915_o_0),
    .B(n_2003_o_0),
    .Y(n_2004_o_0));
 OAI31xp33_ASAP7_75t_R n_2005 (.A1(net8),
    .A2(n_1955_o_0),
    .A3(n_1898_o_0),
    .B(n_2004_o_0),
    .Y(n_2005_o_0));
 NAND3xp33_ASAP7_75t_R n_2006 (.A(n_1936_o_0),
    .B(n_1898_o_0),
    .C(n_1927_o_0),
    .Y(n_2006_o_0));
 INVx1_ASAP7_75t_R n_2007 (.A(n_2006_o_0),
    .Y(n_2007_o_0));
 NOR2xp33_ASAP7_75t_R n_2008 (.A(n_1941_o_0),
    .B(n_1916_o_0),
    .Y(n_2008_o_0));
 NAND2xp33_ASAP7_75t_R n_2009 (.A(n_1916_o_0),
    .B(n_1898_o_0),
    .Y(n_2009_o_0));
 NAND2xp33_ASAP7_75t_R n_2010 (.A(n_1938_o_0),
    .B(n_2009_o_0),
    .Y(n_2010_o_0));
 INVx1_ASAP7_75t_R n_2011 (.A(n_2009_o_0),
    .Y(n_2011_o_0));
 OAI21xp33_ASAP7_75t_R n_2012 (.A1(n_2008_o_0),
    .A2(n_2011_o_0),
    .B(n_1927_o_0),
    .Y(n_2012_o_0));
 OAI211xp5_ASAP7_75t_R n_2013 (.A1(n_2008_o_0),
    .A2(n_2010_o_0),
    .B(n_2012_o_0),
    .C(n_1951_o_0),
    .Y(n_2013_o_0));
 OAI311xp33_ASAP7_75t_R n_2014 (.A1(net98),
    .A2(n_2005_o_0),
    .A3(n_2007_o_0),
    .B1(n_2013_o_0),
    .C1(net31),
    .Y(n_2014_o_0));
 NAND2xp33_ASAP7_75t_R n_2015 (.A(n_1898_o_0),
    .B(n_1938_o_0),
    .Y(n_2015_o_0));
 NOR2xp33_ASAP7_75t_R n_2016 (.A(n_1955_o_0),
    .B(n_2015_o_0),
    .Y(n_2016_o_0));
 NAND2xp33_ASAP7_75t_R n_2017 (.A(n_1890_o_0),
    .B(n_2016_o_0),
    .Y(n_2017_o_0));
 AOI221xp5_ASAP7_75t_R n_2018 (.A1(n_1917_o_0),
    .A2(n_1912_o_0),
    .B1(n_1933_o_0),
    .B2(n_1898_o_0),
    .C(n_1938_o_0),
    .Y(n_2018_o_0));
 NOR3xp33_ASAP7_75t_R n_2019 (.A(n_1937_o_0),
    .B(n_1898_o_0),
    .C(n_1927_o_0),
    .Y(n_2019_o_0));
 OAI221xp5_ASAP7_75t_R n_2020 (.A1(n_1955_o_0),
    .A2(n_2015_o_0),
    .B1(n_2018_o_0),
    .B2(n_2019_o_0),
    .C(n_1890_o_0),
    .Y(n_2020_o_0));
 AOI21xp33_ASAP7_75t_R n_2021 (.A1(n_1895_o_0),
    .A2(n_1897_o_0),
    .B(n_1948_o_0),
    .Y(n_2021_o_0));
 NAND2xp33_ASAP7_75t_R n_2022 (.A(n_1941_o_0),
    .B(n_1932_o_0),
    .Y(n_2022_o_0));
 INVx1_ASAP7_75t_R n_2023 (.A(n_2022_o_0),
    .Y(n_2023_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2024 (.A1(n_1898_o_0),
    .A2(n_1934_o_0),
    .B(net33),
    .C(n_1890_o_0),
    .Y(n_2024_o_0));
 OAI31xp33_ASAP7_75t_R n_2025 (.A1(n_1927_o_0),
    .A2(n_2021_o_0),
    .A3(n_2023_o_0),
    .B(n_2024_o_0),
    .Y(n_2025_o_0));
 AO31x2_ASAP7_75t_R n_2026 (.A1(n_2017_o_0),
    .A2(n_2020_o_0),
    .A3(n_2025_o_0),
    .B(n_1880_o_0),
    .Y(n_2026_o_0));
 INVx1_ASAP7_75t_R n_2027 (.A(n_1865_o_0),
    .Y(n_2027_o_0));
 AOI31xp33_ASAP7_75t_R n_2028 (.A1(n_1872_o_0),
    .A2(n_2014_o_0),
    .A3(n_2026_o_0),
    .B(n_2027_o_0),
    .Y(n_2028_o_0));
 OAI21xp33_ASAP7_75t_R n_2029 (.A1(n_1872_o_0),
    .A2(n_2002_o_0),
    .B(n_2028_o_0),
    .Y(n_2029_o_0));
 OAI21xp33_ASAP7_75t_R n_2030 (.A1(n_1865_o_0),
    .A2(n_1983_o_0),
    .B(n_2029_o_0),
    .Y(n_2030_o_0));
 NOR2xp33_ASAP7_75t_R n_2031 (.A(n_1994_o_0),
    .B(n_1954_o_0),
    .Y(n_2031_o_0));
 AOI31xp33_ASAP7_75t_R n_2032 (.A1(net8),
    .A2(n_2022_o_0),
    .A3(n_2009_o_0),
    .B(n_2031_o_0),
    .Y(n_2032_o_0));
 INVx1_ASAP7_75t_R n_2033 (.A(n_1945_o_0),
    .Y(n_2033_o_0));
 NOR2xp33_ASAP7_75t_R n_2034 (.A(net33),
    .B(n_2033_o_0),
    .Y(n_2034_o_0));
 NAND2xp33_ASAP7_75t_R n_2035 (.A(n_1932_o_0),
    .B(n_1955_o_0),
    .Y(n_2035_o_0));
 NAND2xp33_ASAP7_75t_R n_2036 (.A(n_1927_o_0),
    .B(n_1932_o_0),
    .Y(n_2036_o_0));
 NAND3xp33_ASAP7_75t_R n_2037 (.A(n_1915_o_0),
    .B(n_1898_o_0),
    .C(net33),
    .Y(n_2037_o_0));
 OAI211xp5_ASAP7_75t_R n_2038 (.A1(n_1953_o_0),
    .A2(n_2036_o_0),
    .B(n_1880_o_0),
    .C(n_2037_o_0),
    .Y(n_2038_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2039 (.A1(n_2034_o_0),
    .A2(n_2035_o_0),
    .B(n_2038_o_0),
    .C(net18),
    .Y(n_2039_o_0));
 AOI21xp33_ASAP7_75t_R n_2040 (.A1(n_2032_o_0),
    .A2(n_1993_o_0),
    .B(n_2039_o_0),
    .Y(n_2040_o_0));
 NOR2xp33_ASAP7_75t_R n_2041 (.A(n_1898_o_0),
    .B(n_1927_o_0),
    .Y(n_2041_o_0));
 NOR3xp33_ASAP7_75t_R n_2042 (.A(n_1932_o_0),
    .B(n_1914_o_0),
    .C(n_1927_o_0),
    .Y(n_2042_o_0));
 AOI21xp33_ASAP7_75t_R n_2043 (.A1(n_1936_o_0),
    .A2(n_2041_o_0),
    .B(n_2042_o_0),
    .Y(n_2043_o_0));
 NAND3xp33_ASAP7_75t_R n_2044 (.A(n_1995_o_0),
    .B(n_1993_o_0),
    .C(net33),
    .Y(n_2044_o_0));
 AOI21xp33_ASAP7_75t_R n_2045 (.A1(n_2043_o_0),
    .A2(n_2044_o_0),
    .B(net18),
    .Y(n_2045_o_0));
 NOR3xp33_ASAP7_75t_R n_2046 (.A(n_2040_o_0),
    .B(n_2045_o_0),
    .C(n_1873_o_0),
    .Y(n_2046_o_0));
 OAI21xp33_ASAP7_75t_R n_2047 (.A1(n_1930_o_0),
    .A2(n_1931_o_0),
    .B(n_1934_o_0),
    .Y(n_2047_o_0));
 NAND2xp33_ASAP7_75t_R n_2048 (.A(n_1927_o_0),
    .B(n_2047_o_0),
    .Y(n_2048_o_0));
 NOR2xp33_ASAP7_75t_R n_2049 (.A(n_1898_o_0),
    .B(n_1915_o_0),
    .Y(n_2049_o_0));
 OAI21xp33_ASAP7_75t_R n_2050 (.A1(n_1898_o_0),
    .A2(n_1955_o_0),
    .B(n_1938_o_0),
    .Y(n_2050_o_0));
 NOR2xp33_ASAP7_75t_R n_2051 (.A(n_1914_o_0),
    .B(n_1932_o_0),
    .Y(n_2051_o_0));
 OA21x2_ASAP7_75t_R n_2052 (.A1(n_2050_o_0),
    .A2(n_2051_o_0),
    .B(n_1951_o_0),
    .Y(n_2052_o_0));
 INVx1_ASAP7_75t_R n_2053 (.A(n_1990_o_0),
    .Y(n_2053_o_0));
 NOR4xp25_ASAP7_75t_R n_2054 (.A(n_2053_o_0),
    .B(n_2042_o_0),
    .C(net17),
    .D(n_1918_o_0),
    .Y(n_2054_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2055 (.A1(n_2048_o_0),
    .A2(n_2049_o_0),
    .B(n_2052_o_0),
    .C(n_2054_o_0),
    .Y(n_2055_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2056 (.A1(net8),
    .A2(n_2009_o_0),
    .B(n_2031_o_0),
    .C(n_2035_o_0),
    .Y(n_2056_o_0));
 NOR3xp33_ASAP7_75t_R n_2057 (.A(n_1938_o_0),
    .B(n_1932_o_0),
    .C(n_1955_o_0),
    .Y(n_2057_o_0));
 NAND3xp33_ASAP7_75t_R n_2058 (.A(n_1934_o_0),
    .B(n_1932_o_0),
    .C(n_1927_o_0),
    .Y(n_2058_o_0));
 OAI311xp33_ASAP7_75t_R n_2059 (.A1(n_1898_o_0),
    .A2(net33),
    .A3(n_1917_o_0),
    .B1(n_1951_o_0),
    .C1(n_2058_o_0),
    .Y(n_2059_o_0));
 AOI311xp33_ASAP7_75t_R n_2060 (.A1(net8),
    .A2(n_1955_o_0),
    .A3(n_1898_o_0),
    .B(n_2057_o_0),
    .C(n_2059_o_0),
    .Y(n_2060_o_0));
 AOI211xp5_ASAP7_75t_R n_2061 (.A1(n_2056_o_0),
    .A2(n_1890_o_0),
    .B(n_2060_o_0),
    .C(n_1993_o_0),
    .Y(n_2061_o_0));
 AOI211xp5_ASAP7_75t_R n_2062 (.A1(n_2055_o_0),
    .A2(n_1993_o_0),
    .B(n_1872_o_0),
    .C(n_2061_o_0),
    .Y(n_2062_o_0));
 AOI21xp33_ASAP7_75t_R n_2063 (.A1(n_1938_o_0),
    .A2(n_1918_o_0),
    .B(n_1890_o_0),
    .Y(n_2063_o_0));
 INVx1_ASAP7_75t_R n_2064 (.A(n_2063_o_0),
    .Y(n_2064_o_0));
 NOR2xp33_ASAP7_75t_R n_2065 (.A(n_1898_o_0),
    .B(n_1953_o_0),
    .Y(n_2065_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2066 (.A1(n_1955_o_0),
    .A2(n_2015_o_0),
    .B(n_2048_o_0),
    .C(n_2065_o_0),
    .Y(n_2066_o_0));
 NAND2xp33_ASAP7_75t_R n_2067 (.A(n_1941_o_0),
    .B(n_1916_o_0),
    .Y(n_2067_o_0));
 INVx1_ASAP7_75t_R n_2068 (.A(n_2067_o_0),
    .Y(n_2068_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2069 (.A1(n_2068_o_0),
    .A2(n_2033_o_0),
    .B(net33),
    .C(n_1951_o_0),
    .Y(n_2069_o_0));
 OAI21xp33_ASAP7_75t_R n_2070 (.A1(n_1975_o_0),
    .A2(n_2033_o_0),
    .B(n_2069_o_0),
    .Y(n_2070_o_0));
 OAI21xp33_ASAP7_75t_R n_2071 (.A1(n_2064_o_0),
    .A2(n_2066_o_0),
    .B(n_2070_o_0),
    .Y(n_2071_o_0));
 OAI21xp33_ASAP7_75t_R n_2072 (.A1(n_1898_o_0),
    .A2(n_1934_o_0),
    .B(n_1927_o_0),
    .Y(n_2072_o_0));
 NAND3xp33_ASAP7_75t_R n_2073 (.A(n_1938_o_0),
    .B(n_1898_o_0),
    .C(n_1942_o_0),
    .Y(n_2073_o_0));
 OAI21xp33_ASAP7_75t_R n_2074 (.A1(n_2051_o_0),
    .A2(n_2072_o_0),
    .B(n_2073_o_0),
    .Y(n_2074_o_0));
 NAND2xp33_ASAP7_75t_R n_2075 (.A(n_1912_o_0),
    .B(n_1898_o_0),
    .Y(n_2075_o_0));
 OAI21xp33_ASAP7_75t_R n_2076 (.A1(net4),
    .A2(n_2022_o_0),
    .B(n_1951_o_0),
    .Y(n_2076_o_0));
 INVx1_ASAP7_75t_R n_2077 (.A(n_1943_o_0),
    .Y(n_2077_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2078 (.A1(net4),
    .A2(n_2075_o_0),
    .B(n_2076_o_0),
    .C(n_2077_o_0),
    .Y(n_2078_o_0));
 AOI211xp5_ASAP7_75t_R n_2079 (.A1(n_1890_o_0),
    .A2(n_2074_o_0),
    .B(n_2078_o_0),
    .C(n_1873_o_0),
    .Y(n_2079_o_0));
 AOI21xp33_ASAP7_75t_R n_2080 (.A1(n_1873_o_0),
    .A2(n_2071_o_0),
    .B(n_2079_o_0),
    .Y(n_2080_o_0));
 INVx1_ASAP7_75t_R n_2081 (.A(n_2008_o_0),
    .Y(n_2081_o_0));
 NAND3xp33_ASAP7_75t_R n_2082 (.A(n_2081_o_0),
    .B(n_1949_o_0),
    .C(n_1938_o_0),
    .Y(n_2082_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2083 (.A1(n_1953_o_0),
    .A2(n_2036_o_0),
    .B(n_2082_o_0),
    .C(n_1951_o_0),
    .Y(n_2083_o_0));
 OAI21xp33_ASAP7_75t_R n_2084 (.A1(n_1932_o_0),
    .A2(n_1953_o_0),
    .B(n_1938_o_0),
    .Y(n_2084_o_0));
 INVx1_ASAP7_75t_R n_2085 (.A(n_2084_o_0),
    .Y(n_2085_o_0));
 AOI21xp33_ASAP7_75t_R n_2086 (.A1(n_1978_o_0),
    .A2(n_2085_o_0),
    .B(n_1890_o_0),
    .Y(n_2086_o_0));
 OAI21xp33_ASAP7_75t_R n_2087 (.A1(n_1990_o_0),
    .A2(n_1986_o_0),
    .B(n_2086_o_0),
    .Y(n_2087_o_0));
 OAI21xp33_ASAP7_75t_R n_2088 (.A1(net17),
    .A2(n_2083_o_0),
    .B(n_2087_o_0),
    .Y(n_2088_o_0));
 OAI211xp5_ASAP7_75t_R n_2089 (.A1(n_1898_o_0),
    .A2(n_1915_o_0),
    .B(n_2047_o_0),
    .C(n_1927_o_0),
    .Y(n_2089_o_0));
 OAI31xp33_ASAP7_75t_R n_2090 (.A1(net33),
    .A2(n_1932_o_0),
    .A3(n_1942_o_0),
    .B(n_2089_o_0),
    .Y(n_2090_o_0));
 OAI211xp5_ASAP7_75t_R n_2091 (.A1(n_1898_o_0),
    .A2(n_1916_o_0),
    .B(n_1927_o_0),
    .C(n_1941_o_0),
    .Y(n_2091_o_0));
 OAI211xp5_ASAP7_75t_R n_2092 (.A1(n_2015_o_0),
    .A2(n_1914_o_0),
    .B(n_2091_o_0),
    .C(n_1951_o_0),
    .Y(n_2092_o_0));
 OAI211xp5_ASAP7_75t_R n_2093 (.A1(n_2090_o_0),
    .A2(n_1951_o_0),
    .B(n_2092_o_0),
    .C(n_1873_o_0),
    .Y(n_2093_o_0));
 OAI211xp5_ASAP7_75t_R n_2094 (.A1(n_2088_o_0),
    .A2(n_1873_o_0),
    .B(net31),
    .C(n_2093_o_0),
    .Y(n_2094_o_0));
 OAI211xp5_ASAP7_75t_R n_2095 (.A1(net31),
    .A2(n_2080_o_0),
    .B(n_2094_o_0),
    .C(n_2027_o_0),
    .Y(n_2095_o_0));
 OAI31xp33_ASAP7_75t_R n_2096 (.A1(n_2027_o_0),
    .A2(n_2046_o_0),
    .A3(n_2062_o_0),
    .B(n_2095_o_0),
    .Y(n_2096_o_0));
 INVx1_ASAP7_75t_R n_2097 (.A(n_2035_o_0),
    .Y(n_2097_o_0));
 NAND2xp33_ASAP7_75t_R n_2098 (.A(n_1938_o_0),
    .B(n_1998_o_0),
    .Y(n_2098_o_0));
 OAI211xp5_ASAP7_75t_R n_2099 (.A1(n_2097_o_0),
    .A2(n_2098_o_0),
    .B(n_2058_o_0),
    .C(n_1951_o_0),
    .Y(n_2099_o_0));
 NAND3xp33_ASAP7_75t_R n_2100 (.A(n_2081_o_0),
    .B(n_1949_o_0),
    .C(net33),
    .Y(n_2100_o_0));
 OAI21xp33_ASAP7_75t_R n_2101 (.A1(net33),
    .A2(n_1994_o_0),
    .B(n_2100_o_0),
    .Y(n_2101_o_0));
 OAI22xp33_ASAP7_75t_R n_2102 (.A1(n_2099_o_0),
    .A2(n_2007_o_0),
    .B1(n_2101_o_0),
    .B2(net98),
    .Y(n_2102_o_0));
 NOR2xp33_ASAP7_75t_R n_2103 (.A(n_1942_o_0),
    .B(n_1932_o_0),
    .Y(n_2103_o_0));
 OAI22xp33_ASAP7_75t_R n_2104 (.A1(n_2072_o_0),
    .A2(n_2103_o_0),
    .B1(n_1949_o_0),
    .B2(net33),
    .Y(n_2104_o_0));
 AO21x1_ASAP7_75t_R n_2105 (.A1(n_2022_o_0),
    .A2(n_2009_o_0),
    .B(n_1938_o_0),
    .Y(n_2105_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2106 (.A1(n_2105_o_0),
    .A2(n_1950_o_0),
    .B(n_1890_o_0),
    .C(n_1880_o_0),
    .Y(n_2106_o_0));
 AOI21xp33_ASAP7_75t_R n_2107 (.A1(n_2104_o_0),
    .A2(n_1890_o_0),
    .B(n_2106_o_0),
    .Y(n_2107_o_0));
 AOI21xp33_ASAP7_75t_R n_2108 (.A1(n_1993_o_0),
    .A2(n_2102_o_0),
    .B(n_2107_o_0),
    .Y(n_2108_o_0));
 INVx1_ASAP7_75t_R n_2109 (.A(n_1935_o_0),
    .Y(n_2109_o_0));
 AOI21xp33_ASAP7_75t_R n_2110 (.A1(n_1916_o_0),
    .A2(n_1912_o_0),
    .B(n_1898_o_0),
    .Y(n_2110_o_0));
 OAI21xp33_ASAP7_75t_R n_2111 (.A1(n_1916_o_0),
    .A2(n_1932_o_0),
    .B(n_1938_o_0),
    .Y(n_2111_o_0));
 NOR2xp33_ASAP7_75t_R n_2112 (.A(n_2110_o_0),
    .B(n_2111_o_0),
    .Y(n_2112_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2113 (.A1(n_1898_o_0),
    .A2(n_1948_o_0),
    .B(n_2109_o_0),
    .C(n_2112_o_0),
    .Y(n_2113_o_0));
 OAI21xp33_ASAP7_75t_R n_2114 (.A1(n_1932_o_0),
    .A2(n_1936_o_0),
    .B(net33),
    .Y(n_2114_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2115 (.A1(n_1912_o_0),
    .A2(n_1932_o_0),
    .B(n_1917_o_0),
    .C(n_1938_o_0),
    .D(n_1890_o_0),
    .Y(n_2115_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2116 (.A1(n_1994_o_0),
    .A2(n_2114_o_0),
    .B(n_2115_o_0),
    .C(n_1993_o_0),
    .Y(n_2116_o_0));
 OAI21xp33_ASAP7_75t_R n_2117 (.A1(net98),
    .A2(n_2113_o_0),
    .B(n_2116_o_0),
    .Y(n_2117_o_0));
 AOI211xp5_ASAP7_75t_R n_2118 (.A1(n_1916_o_0),
    .A2(n_1932_o_0),
    .B(n_1938_o_0),
    .C(n_1912_o_0),
    .Y(n_2118_o_0));
 NOR2xp33_ASAP7_75t_R n_2119 (.A(n_1898_o_0),
    .B(n_1927_o_0),
    .Y(n_2119_o_0));
 AOI21xp33_ASAP7_75t_R n_2120 (.A1(n_1914_o_0),
    .A2(n_2119_o_0),
    .B(n_1890_o_0),
    .Y(n_2120_o_0));
 OAI31xp33_ASAP7_75t_R n_2121 (.A1(n_1938_o_0),
    .A2(n_2033_o_0),
    .A3(n_2065_o_0),
    .B(n_2120_o_0),
    .Y(n_2121_o_0));
 OAI31xp33_ASAP7_75t_R n_2122 (.A1(n_1951_o_0),
    .A2(n_1943_o_0),
    .A3(n_2118_o_0),
    .B(n_2121_o_0),
    .Y(n_2122_o_0));
 OAI311xp33_ASAP7_75t_R n_2123 (.A1(n_1936_o_0),
    .A2(n_1932_o_0),
    .A3(net33),
    .B1(n_1993_o_0),
    .C1(n_2122_o_0),
    .Y(n_2123_o_0));
 AO21x1_ASAP7_75t_R n_2124 (.A1(n_2117_o_0),
    .A2(n_2123_o_0),
    .B(n_2027_o_0),
    .Y(n_2124_o_0));
 OAI21xp33_ASAP7_75t_R n_2125 (.A1(n_1865_o_0),
    .A2(n_2108_o_0),
    .B(n_2124_o_0),
    .Y(n_2125_o_0));
 OAI21xp33_ASAP7_75t_R n_2126 (.A1(n_1898_o_0),
    .A2(n_1942_o_0),
    .B(n_1938_o_0),
    .Y(n_2126_o_0));
 OAI21xp33_ASAP7_75t_R n_2127 (.A1(net8),
    .A2(n_1973_o_0),
    .B(n_2126_o_0),
    .Y(n_2127_o_0));
 AOI31xp33_ASAP7_75t_R n_2128 (.A1(n_1927_o_0),
    .A2(n_1984_o_0),
    .A3(n_1949_o_0),
    .B(n_1890_o_0),
    .Y(n_2128_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2129 (.A1(n_2022_o_0),
    .A2(net33),
    .B(n_2128_o_0),
    .C(n_1880_o_0),
    .Y(n_2129_o_0));
 OAI21xp33_ASAP7_75t_R n_2130 (.A1(n_2127_o_0),
    .A2(net18),
    .B(n_2129_o_0),
    .Y(n_2130_o_0));
 OAI22xp33_ASAP7_75t_R n_2131 (.A1(n_1990_o_0),
    .A2(n_2065_o_0),
    .B1(n_2015_o_0),
    .B2(n_1955_o_0),
    .Y(n_2131_o_0));
 OAI21xp33_ASAP7_75t_R n_2132 (.A1(n_1898_o_0),
    .A2(n_1915_o_0),
    .B(n_1927_o_0),
    .Y(n_2132_o_0));
 AOI211xp5_ASAP7_75t_R n_2133 (.A1(n_2041_o_0),
    .A2(n_1936_o_0),
    .B(n_2042_o_0),
    .C(n_1890_o_0),
    .Y(n_2133_o_0));
 OAI21xp33_ASAP7_75t_R n_2134 (.A1(n_2132_o_0),
    .A2(n_2011_o_0),
    .B(n_2133_o_0),
    .Y(n_2134_o_0));
 OAI211xp5_ASAP7_75t_R n_2135 (.A1(n_2131_o_0),
    .A2(net17),
    .B(n_2134_o_0),
    .C(net31),
    .Y(n_2135_o_0));
 NAND3xp33_ASAP7_75t_R n_2136 (.A(n_2130_o_0),
    .B(n_2135_o_0),
    .C(n_2027_o_0),
    .Y(n_2136_o_0));
 AOI21xp33_ASAP7_75t_R n_2137 (.A1(n_1915_o_0),
    .A2(n_1932_o_0),
    .B(n_2084_o_0),
    .Y(n_2137_o_0));
 AOI31xp33_ASAP7_75t_R n_2138 (.A1(n_1949_o_0),
    .A2(n_1984_o_0),
    .A3(net33),
    .B(n_2137_o_0),
    .Y(n_2138_o_0));
 OAI21xp33_ASAP7_75t_R n_2139 (.A1(n_2103_o_0),
    .A2(n_2065_o_0),
    .B(n_1927_o_0),
    .Y(n_2139_o_0));
 AOI31xp33_ASAP7_75t_R n_2140 (.A1(n_1890_o_0),
    .A2(n_2139_o_0),
    .A3(n_1950_o_0),
    .B(n_1880_o_0),
    .Y(n_2140_o_0));
 OAI21xp33_ASAP7_75t_R n_2141 (.A1(n_1890_o_0),
    .A2(n_2138_o_0),
    .B(n_2140_o_0),
    .Y(n_2141_o_0));
 NAND2xp33_ASAP7_75t_R n_2142 (.A(n_1927_o_0),
    .B(n_2009_o_0),
    .Y(n_2142_o_0));
 AOI21xp33_ASAP7_75t_R n_2143 (.A1(n_1932_o_0),
    .A2(n_1955_o_0),
    .B(n_2142_o_0),
    .Y(n_2143_o_0));
 OAI31xp33_ASAP7_75t_R n_2144 (.A1(net33),
    .A2(n_2021_o_0),
    .A3(n_1994_o_0),
    .B(net17),
    .Y(n_2144_o_0));
 OAI21xp33_ASAP7_75t_R n_2145 (.A1(n_2051_o_0),
    .A2(n_2132_o_0),
    .B(n_2126_o_0),
    .Y(n_2145_o_0));
 AOI21xp33_ASAP7_75t_R n_2146 (.A1(n_1890_o_0),
    .A2(n_2145_o_0),
    .B(n_1993_o_0),
    .Y(n_2146_o_0));
 OAI21xp33_ASAP7_75t_R n_2147 (.A1(n_2143_o_0),
    .A2(n_2144_o_0),
    .B(n_2146_o_0),
    .Y(n_2147_o_0));
 AO21x1_ASAP7_75t_R n_2148 (.A1(n_2141_o_0),
    .A2(n_2147_o_0),
    .B(n_2027_o_0),
    .Y(n_2148_o_0));
 AOI21xp33_ASAP7_75t_R n_2149 (.A1(n_2136_o_0),
    .A2(n_2148_o_0),
    .B(n_1873_o_0),
    .Y(n_2149_o_0));
 AOI21xp33_ASAP7_75t_R n_2150 (.A1(n_1873_o_0),
    .A2(n_2125_o_0),
    .B(n_2149_o_0),
    .Y(n_2150_o_0));
 OAI21xp33_ASAP7_75t_R n_2151 (.A1(n_2008_o_0),
    .A2(n_1918_o_0),
    .B(n_1938_o_0),
    .Y(n_2151_o_0));
 OA211x2_ASAP7_75t_R n_2152 (.A1(n_1990_o_0),
    .A2(n_1994_o_0),
    .B(n_2151_o_0),
    .C(n_1890_o_0),
    .Y(n_2152_o_0));
 INVx1_ASAP7_75t_R n_2153 (.A(n_2072_o_0),
    .Y(n_2153_o_0));
 AOI21xp33_ASAP7_75t_R n_2154 (.A1(n_2009_o_0),
    .A2(n_2022_o_0),
    .B(net33),
    .Y(n_2154_o_0));
 NOR3xp33_ASAP7_75t_R n_2155 (.A(n_2153_o_0),
    .B(n_1890_o_0),
    .C(n_2154_o_0),
    .Y(n_2155_o_0));
 OAI22xp33_ASAP7_75t_R n_2156 (.A1(n_2015_o_0),
    .A2(n_1937_o_0),
    .B1(n_2036_o_0),
    .B2(n_1934_o_0),
    .Y(n_2156_o_0));
 NAND3xp33_ASAP7_75t_R n_2157 (.A(n_2047_o_0),
    .B(n_1995_o_0),
    .C(n_1938_o_0),
    .Y(n_2157_o_0));
 OAI31xp33_ASAP7_75t_R n_2158 (.A1(n_2051_o_0),
    .A2(n_2065_o_0),
    .A3(net8),
    .B(n_2157_o_0),
    .Y(n_2158_o_0));
 OAI321xp33_ASAP7_75t_R n_2159 (.A1(n_2156_o_0),
    .A2(n_2057_o_0),
    .A3(n_2064_o_0),
    .B1(n_2158_o_0),
    .B2(n_1951_o_0),
    .C(n_1880_o_0),
    .Y(n_2159_o_0));
 OAI31xp33_ASAP7_75t_R n_2160 (.A1(net31),
    .A2(n_2152_o_0),
    .A3(n_2155_o_0),
    .B(n_2159_o_0),
    .Y(n_2160_o_0));
 INVx1_ASAP7_75t_R n_2161 (.A(n_1968_o_0),
    .Y(n_2161_o_0));
 OAI31xp33_ASAP7_75t_R n_2162 (.A1(net33),
    .A2(n_2021_o_0),
    .A3(n_2161_o_0),
    .B(n_1951_o_0),
    .Y(n_2162_o_0));
 INVx1_ASAP7_75t_R n_2163 (.A(n_2091_o_0),
    .Y(n_2163_o_0));
 INVx1_ASAP7_75t_R n_2164 (.A(n_1984_o_0),
    .Y(n_2164_o_0));
 OAI21xp33_ASAP7_75t_R n_2165 (.A1(net8),
    .A2(n_2164_o_0),
    .B(n_2151_o_0),
    .Y(n_2165_o_0));
 OAI22xp33_ASAP7_75t_R n_2166 (.A1(n_2162_o_0),
    .A2(n_2163_o_0),
    .B1(n_2165_o_0),
    .B2(n_1951_o_0),
    .Y(n_2166_o_0));
 OAI21xp33_ASAP7_75t_R n_2167 (.A1(n_1932_o_0),
    .A2(n_1934_o_0),
    .B(n_1938_o_0),
    .Y(n_2167_o_0));
 INVx1_ASAP7_75t_R n_2168 (.A(n_2167_o_0),
    .Y(n_2168_o_0));
 OAI21xp33_ASAP7_75t_R n_2169 (.A1(n_1898_o_0),
    .A2(n_1937_o_0),
    .B(n_2168_o_0),
    .Y(n_2169_o_0));
 AOI21xp33_ASAP7_75t_R n_2170 (.A1(n_1941_o_0),
    .A2(n_1917_o_0),
    .B(n_1898_o_0),
    .Y(n_2170_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2171 (.A1(n_2170_o_0),
    .A2(net4),
    .B(n_1975_o_0),
    .C(n_2042_o_0),
    .Y(n_2171_o_0));
 NOR2xp33_ASAP7_75t_R n_2172 (.A(n_1890_o_0),
    .B(n_1993_o_0),
    .Y(n_2172_o_0));
 AOI31xp33_ASAP7_75t_R n_2173 (.A1(n_2006_o_0),
    .A2(n_2171_o_0),
    .A3(net31),
    .B(n_2172_o_0),
    .Y(n_2173_o_0));
 AOI31xp33_ASAP7_75t_R n_2174 (.A1(n_2012_o_0),
    .A2(n_2169_o_0),
    .A3(net98),
    .B(n_2173_o_0),
    .Y(n_2174_o_0));
 AOI211xp5_ASAP7_75t_R n_2175 (.A1(n_2166_o_0),
    .A2(n_1993_o_0),
    .B(n_2174_o_0),
    .C(n_1872_o_0),
    .Y(n_2175_o_0));
 AOI21xp33_ASAP7_75t_R n_2176 (.A1(n_1872_o_0),
    .A2(n_2160_o_0),
    .B(n_2175_o_0),
    .Y(n_2176_o_0));
 INVx1_ASAP7_75t_R n_2177 (.A(n_2115_o_0),
    .Y(n_2177_o_0));
 OAI211xp5_ASAP7_75t_R n_2178 (.A1(n_1937_o_0),
    .A2(n_1898_o_0),
    .B(n_2009_o_0),
    .C(n_1927_o_0),
    .Y(n_2178_o_0));
 AO21x1_ASAP7_75t_R n_2179 (.A1(n_2178_o_0),
    .A2(n_2043_o_0),
    .B(net98),
    .Y(n_2179_o_0));
 AOI21xp33_ASAP7_75t_R n_2180 (.A1(n_2082_o_0),
    .A2(n_1977_o_0),
    .B(n_1951_o_0),
    .Y(n_2180_o_0));
 OAI21xp33_ASAP7_75t_R n_2181 (.A1(n_1932_o_0),
    .A2(n_1934_o_0),
    .B(n_1938_o_0),
    .Y(n_2181_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2182 (.A1(n_1937_o_0),
    .A2(n_1898_o_0),
    .B(n_1986_o_0),
    .C(n_1927_o_0),
    .Y(n_2182_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2183 (.A1(n_1989_o_0),
    .A2(n_2181_o_0),
    .B(n_2182_o_0),
    .C(n_1890_o_0),
    .Y(n_2183_o_0));
 NOR3xp33_ASAP7_75t_R n_2184 (.A(n_2180_o_0),
    .B(n_2183_o_0),
    .C(n_1993_o_0),
    .Y(n_2184_o_0));
 AOI31xp33_ASAP7_75t_R n_2185 (.A1(n_1993_o_0),
    .A2(n_2177_o_0),
    .A3(n_2179_o_0),
    .B(n_2184_o_0),
    .Y(n_2185_o_0));
 NOR3xp33_ASAP7_75t_R n_2186 (.A(n_1938_o_0),
    .B(n_1936_o_0),
    .C(n_1932_o_0),
    .Y(n_2186_o_0));
 OAI221xp5_ASAP7_75t_R n_2187 (.A1(n_1989_o_0),
    .A2(n_2142_o_0),
    .B1(n_1986_o_0),
    .B2(n_2181_o_0),
    .C(n_1993_o_0),
    .Y(n_2187_o_0));
 OAI31xp33_ASAP7_75t_R n_2188 (.A1(n_2112_o_0),
    .A2(n_2186_o_0),
    .A3(n_1993_o_0),
    .B(n_2187_o_0),
    .Y(n_2188_o_0));
 NOR3xp33_ASAP7_75t_R n_2189 (.A(n_1934_o_0),
    .B(n_1932_o_0),
    .C(n_1927_o_0),
    .Y(n_2189_o_0));
 OAI22xp33_ASAP7_75t_R n_2190 (.A1(n_1973_o_0),
    .A2(n_1963_o_0),
    .B1(n_2036_o_0),
    .B2(n_1934_o_0),
    .Y(n_2190_o_0));
 AO21x1_ASAP7_75t_R n_2191 (.A1(n_2190_o_0),
    .A2(n_1993_o_0),
    .B(n_1966_o_0),
    .Y(n_2191_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2192 (.A1(n_1880_o_0),
    .A2(n_2189_o_0),
    .B(n_2191_o_0),
    .C(net17),
    .Y(n_2192_o_0));
 OAI211xp5_ASAP7_75t_R n_2193 (.A1(n_2188_o_0),
    .A2(net98),
    .B(n_2192_o_0),
    .C(n_1872_o_0),
    .Y(n_2193_o_0));
 OAI211xp5_ASAP7_75t_R n_2194 (.A1(n_2185_o_0),
    .A2(n_1872_o_0),
    .B(n_1865_o_0),
    .C(n_2193_o_0),
    .Y(n_2194_o_0));
 OAI21xp33_ASAP7_75t_R n_2195 (.A1(n_1865_o_0),
    .A2(n_2176_o_0),
    .B(n_2194_o_0),
    .Y(n_2195_o_0));
 OAI21xp33_ASAP7_75t_R n_2196 (.A1(n_1932_o_0),
    .A2(n_1953_o_0),
    .B(n_1938_o_0),
    .Y(n_2196_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2197 (.A1(n_1932_o_0),
    .A2(n_1934_o_0),
    .B(n_2196_o_0),
    .C(n_1928_o_0),
    .Y(n_2197_o_0));
 OA21x2_ASAP7_75t_R n_2198 (.A1(n_2010_o_0),
    .A2(n_1989_o_0),
    .B(n_1993_o_0),
    .Y(n_2198_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2199 (.A1(net8),
    .A2(n_1898_o_0),
    .B(n_2198_o_0),
    .C(net98),
    .Y(n_2199_o_0));
 NOR3xp33_ASAP7_75t_R n_2200 (.A(n_1927_o_0),
    .B(n_1898_o_0),
    .C(n_1941_o_0),
    .Y(n_2200_o_0));
 NOR4xp25_ASAP7_75t_R n_2201 (.A(n_2016_o_0),
    .B(n_2031_o_0),
    .C(n_2200_o_0),
    .D(n_1880_o_0),
    .Y(n_2201_o_0));
 AOI311xp33_ASAP7_75t_R n_2202 (.A1(net31),
    .A2(n_2050_o_0),
    .A3(n_2132_o_0),
    .B(n_1890_o_0),
    .C(n_2201_o_0),
    .Y(n_2202_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2203 (.A1(n_1993_o_0),
    .A2(n_2197_o_0),
    .B(n_2199_o_0),
    .C(n_2202_o_0),
    .Y(n_2203_o_0));
 AO21x1_ASAP7_75t_R n_2204 (.A1(n_1957_o_0),
    .A2(n_2012_o_0),
    .B(net31),
    .Y(n_2204_o_0));
 OAI211xp5_ASAP7_75t_R n_2205 (.A1(net33),
    .A2(n_1915_o_0),
    .B(n_2058_o_0),
    .C(net31),
    .Y(n_2205_o_0));
 INVx1_ASAP7_75t_R n_2206 (.A(n_2178_o_0),
    .Y(n_2206_o_0));
 AOI21xp33_ASAP7_75t_R n_2207 (.A1(n_2067_o_0),
    .A2(n_1998_o_0),
    .B(n_1927_o_0),
    .Y(n_2207_o_0));
 OAI211xp5_ASAP7_75t_R n_2208 (.A1(n_1937_o_0),
    .A2(n_1898_o_0),
    .B(n_2075_o_0),
    .C(n_1927_o_0),
    .Y(n_2208_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2209 (.A1(n_2208_o_0),
    .A2(n_2073_o_0),
    .B(n_1993_o_0),
    .C(n_1951_o_0),
    .Y(n_2209_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2210 (.A1(n_2206_o_0),
    .A2(n_2207_o_0),
    .B(n_1993_o_0),
    .C(n_2209_o_0),
    .Y(n_2210_o_0));
 AOI31xp33_ASAP7_75t_R n_2211 (.A1(n_1890_o_0),
    .A2(n_2204_o_0),
    .A3(n_2205_o_0),
    .B(n_2210_o_0),
    .Y(n_2211_o_0));
 OAI21xp33_ASAP7_75t_R n_2212 (.A1(n_1873_o_0),
    .A2(n_2211_o_0),
    .B(n_1865_o_0),
    .Y(n_2212_o_0));
 OAI211xp5_ASAP7_75t_R n_2213 (.A1(net4),
    .A2(n_2022_o_0),
    .B(n_2073_o_0),
    .C(n_1890_o_0),
    .Y(n_2213_o_0));
 NOR2xp33_ASAP7_75t_R n_2214 (.A(n_2057_o_0),
    .B(n_2213_o_0),
    .Y(n_2214_o_0));
 NAND2xp33_ASAP7_75t_R n_2215 (.A(n_1927_o_0),
    .B(n_1962_o_0),
    .Y(n_2215_o_0));
 INVx1_ASAP7_75t_R n_2216 (.A(n_2215_o_0),
    .Y(n_2216_o_0));
 OAI21xp33_ASAP7_75t_R n_2217 (.A1(n_1989_o_0),
    .A2(n_2084_o_0),
    .B(n_1951_o_0),
    .Y(n_2217_o_0));
 AOI21xp33_ASAP7_75t_R n_2218 (.A1(n_1995_o_0),
    .A2(n_2216_o_0),
    .B(n_2217_o_0),
    .Y(n_2218_o_0));
 AOI211xp5_ASAP7_75t_R n_2219 (.A1(n_2214_o_0),
    .A2(n_2077_o_0),
    .B(net31),
    .C(n_2218_o_0),
    .Y(n_2219_o_0));
 OAI21xp33_ASAP7_75t_R n_2220 (.A1(n_1932_o_0),
    .A2(n_1914_o_0),
    .B(n_1938_o_0),
    .Y(n_2220_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2221 (.A1(n_1948_o_0),
    .A2(n_1932_o_0),
    .B(n_2220_o_0),
    .C(n_1969_o_0),
    .Y(n_2221_o_0));
 OAI211xp5_ASAP7_75t_R n_2222 (.A1(n_1932_o_0),
    .A2(n_1936_o_0),
    .B(n_2077_o_0),
    .C(n_1951_o_0),
    .Y(n_2222_o_0));
 INVx1_ASAP7_75t_R n_2223 (.A(n_2058_o_0),
    .Y(n_2223_o_0));
 OAI22xp33_ASAP7_75t_R n_2224 (.A1(n_2221_o_0),
    .A2(n_1951_o_0),
    .B1(n_2222_o_0),
    .B2(n_2223_o_0),
    .Y(n_2224_o_0));
 OAI21xp33_ASAP7_75t_R n_2225 (.A1(n_1993_o_0),
    .A2(n_2224_o_0),
    .B(n_1872_o_0),
    .Y(n_2225_o_0));
 AOI21xp33_ASAP7_75t_R n_2226 (.A1(n_1927_o_0),
    .A2(n_1968_o_0),
    .B(n_1890_o_0),
    .Y(n_2226_o_0));
 OAI21xp33_ASAP7_75t_R n_2227 (.A1(n_1965_o_0),
    .A2(n_1932_o_0),
    .B(n_2226_o_0),
    .Y(n_2227_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2228 (.A1(n_1994_o_0),
    .A2(n_2011_o_0),
    .B(net33),
    .C(n_1951_o_0),
    .Y(n_2228_o_0));
 OAI31xp33_ASAP7_75t_R n_2229 (.A1(net33),
    .A2(n_2033_o_0),
    .A3(n_2097_o_0),
    .B(n_2228_o_0),
    .Y(n_2229_o_0));
 AOI21xp33_ASAP7_75t_R n_2230 (.A1(n_2227_o_0),
    .A2(n_2229_o_0),
    .B(n_1993_o_0),
    .Y(n_2230_o_0));
 NAND3xp33_ASAP7_75t_R n_2231 (.A(n_2022_o_0),
    .B(n_2009_o_0),
    .C(n_1938_o_0),
    .Y(n_2231_o_0));
 OAI31xp33_ASAP7_75t_R n_2232 (.A1(n_1973_o_0),
    .A2(n_2008_o_0),
    .A3(net8),
    .B(n_2231_o_0),
    .Y(n_2232_o_0));
 OAI31xp33_ASAP7_75t_R n_2233 (.A1(net4),
    .A2(n_1973_o_0),
    .A3(n_1956_o_0),
    .B(n_1951_o_0),
    .Y(n_2233_o_0));
 OAI21xp33_ASAP7_75t_R n_2234 (.A1(n_2207_o_0),
    .A2(n_2233_o_0),
    .B(n_1993_o_0),
    .Y(n_2234_o_0));
 AOI21xp33_ASAP7_75t_R n_2235 (.A1(n_1890_o_0),
    .A2(n_2232_o_0),
    .B(n_2234_o_0),
    .Y(n_2235_o_0));
 OAI21xp33_ASAP7_75t_R n_2236 (.A1(n_2230_o_0),
    .A2(n_2235_o_0),
    .B(n_1873_o_0),
    .Y(n_2236_o_0));
 OAI211xp5_ASAP7_75t_R n_2237 (.A1(n_2219_o_0),
    .A2(n_2225_o_0),
    .B(n_2236_o_0),
    .C(n_2027_o_0),
    .Y(n_2237_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2238 (.A1(n_1873_o_0),
    .A2(n_2203_o_0),
    .B(n_2212_o_0),
    .C(n_2237_o_0),
    .Y(n_2238_o_0));
 NOR2xp33_ASAP7_75t_R n_2239 (.A(n_1927_o_0),
    .B(n_1986_o_0),
    .Y(n_2239_o_0));
 OAI21xp33_ASAP7_75t_R n_2240 (.A1(n_1914_o_0),
    .A2(n_1932_o_0),
    .B(n_1927_o_0),
    .Y(n_2240_o_0));
 AOI21xp33_ASAP7_75t_R n_2241 (.A1(n_1932_o_0),
    .A2(n_1936_o_0),
    .B(n_2240_o_0),
    .Y(n_2241_o_0));
 AOI21xp33_ASAP7_75t_R n_2242 (.A1(n_2239_o_0),
    .A2(n_2067_o_0),
    .B(n_2241_o_0),
    .Y(n_2242_o_0));
 NOR2xp33_ASAP7_75t_R n_2243 (.A(n_2110_o_0),
    .B(n_2103_o_0),
    .Y(n_2243_o_0));
 AOI21xp33_ASAP7_75t_R n_2244 (.A1(n_2243_o_0),
    .A2(net4),
    .B(n_1872_o_0),
    .Y(n_2244_o_0));
 OAI21xp33_ASAP7_75t_R n_2245 (.A1(n_2142_o_0),
    .A2(n_2065_o_0),
    .B(n_2244_o_0),
    .Y(n_2245_o_0));
 OAI21xp33_ASAP7_75t_R n_2246 (.A1(n_1873_o_0),
    .A2(n_2242_o_0),
    .B(n_2245_o_0),
    .Y(n_2246_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2247 (.A1(net8),
    .A2(n_1916_o_0),
    .B(n_1912_o_0),
    .C(n_1872_o_0),
    .Y(n_2247_o_0));
 OAI211xp5_ASAP7_75t_R n_2248 (.A1(n_1989_o_0),
    .A2(n_1954_o_0),
    .B(n_1873_o_0),
    .C(n_1970_o_0),
    .Y(n_2248_o_0));
 OAI21xp33_ASAP7_75t_R n_2249 (.A1(net33),
    .A2(n_1995_o_0),
    .B(n_1890_o_0),
    .Y(n_2249_o_0));
 AOI21xp33_ASAP7_75t_R n_2250 (.A1(n_2247_o_0),
    .A2(n_2248_o_0),
    .B(n_2249_o_0),
    .Y(n_2250_o_0));
 AOI21xp33_ASAP7_75t_R n_2251 (.A1(net18),
    .A2(n_2246_o_0),
    .B(n_2250_o_0),
    .Y(n_2251_o_0));
 INVx1_ASAP7_75t_R n_2252 (.A(n_2142_o_0),
    .Y(n_2252_o_0));
 OAI21xp33_ASAP7_75t_R n_2253 (.A1(n_1914_o_0),
    .A2(n_2015_o_0),
    .B(n_1890_o_0),
    .Y(n_2253_o_0));
 OAI211xp5_ASAP7_75t_R n_2254 (.A1(n_1989_o_0),
    .A2(net4),
    .B(n_2077_o_0),
    .C(n_1951_o_0),
    .Y(n_2254_o_0));
 OAI31xp33_ASAP7_75t_R n_2255 (.A1(n_2252_o_0),
    .A2(n_2170_o_0),
    .A3(n_2253_o_0),
    .B(n_2254_o_0),
    .Y(n_2255_o_0));
 AOI31xp33_ASAP7_75t_R n_2256 (.A1(net8),
    .A2(n_1968_o_0),
    .A3(n_1998_o_0),
    .B(n_1890_o_0),
    .Y(n_2256_o_0));
 OAI21xp33_ASAP7_75t_R n_2257 (.A1(n_2164_o_0),
    .A2(n_1990_o_0),
    .B(n_2256_o_0),
    .Y(n_2257_o_0));
 OAI21xp33_ASAP7_75t_R n_2258 (.A1(n_2008_o_0),
    .A2(n_2010_o_0),
    .B(n_1890_o_0),
    .Y(n_2258_o_0));
 AO21x1_ASAP7_75t_R n_2259 (.A1(net33),
    .A2(n_1916_o_0),
    .B(n_2258_o_0),
    .Y(n_2259_o_0));
 AOI31xp33_ASAP7_75t_R n_2260 (.A1(n_2257_o_0),
    .A2(n_2259_o_0),
    .A3(n_1873_o_0),
    .B(n_2027_o_0),
    .Y(n_2260_o_0));
 OAI21xp33_ASAP7_75t_R n_2261 (.A1(n_2255_o_0),
    .A2(n_1873_o_0),
    .B(n_2260_o_0),
    .Y(n_2261_o_0));
 OAI21xp33_ASAP7_75t_R n_2262 (.A1(n_1865_o_0),
    .A2(n_2251_o_0),
    .B(n_2261_o_0),
    .Y(n_2262_o_0));
 NOR2xp33_ASAP7_75t_R n_2263 (.A(n_2050_o_0),
    .B(n_1973_o_0),
    .Y(n_2263_o_0));
 OAI321xp33_ASAP7_75t_R n_2264 (.A1(n_1898_o_0),
    .A2(n_1915_o_0),
    .A3(net33),
    .B1(n_2048_o_0),
    .B2(n_2097_o_0),
    .C(n_1890_o_0),
    .Y(n_2264_o_0));
 OAI31xp33_ASAP7_75t_R n_2265 (.A1(n_2223_o_0),
    .A2(n_2263_o_0),
    .A3(n_1890_o_0),
    .B(n_2264_o_0),
    .Y(n_2265_o_0));
 NAND3xp33_ASAP7_75t_R n_2266 (.A(n_2167_o_0),
    .B(n_2182_o_0),
    .C(n_1890_o_0),
    .Y(n_2266_o_0));
 OAI211xp5_ASAP7_75t_R n_2267 (.A1(n_1953_o_0),
    .A2(n_1898_o_0),
    .B(n_2196_o_0),
    .C(n_1951_o_0),
    .Y(n_2267_o_0));
 AOI31xp33_ASAP7_75t_R n_2268 (.A1(n_1873_o_0),
    .A2(n_2266_o_0),
    .A3(n_2267_o_0),
    .B(n_1865_o_0),
    .Y(n_2268_o_0));
 OAI21xp33_ASAP7_75t_R n_2269 (.A1(n_2265_o_0),
    .A2(n_1873_o_0),
    .B(n_2268_o_0),
    .Y(n_2269_o_0));
 AOI21xp33_ASAP7_75t_R n_2270 (.A1(n_1932_o_0),
    .A2(n_1937_o_0),
    .B(n_1990_o_0),
    .Y(n_2270_o_0));
 INVx1_ASAP7_75t_R n_2271 (.A(n_2120_o_0),
    .Y(n_2271_o_0));
 NOR3xp33_ASAP7_75t_R n_2272 (.A(n_1915_o_0),
    .B(n_1932_o_0),
    .C(n_1927_o_0),
    .Y(n_2272_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2273 (.A1(net33),
    .A2(n_1937_o_0),
    .B(n_2272_o_0),
    .C(n_1890_o_0),
    .Y(n_2273_o_0));
 OAI31xp33_ASAP7_75t_R n_2274 (.A1(n_2189_o_0),
    .A2(n_2270_o_0),
    .A3(n_2271_o_0),
    .B(n_2273_o_0),
    .Y(n_2274_o_0));
 OAI21xp33_ASAP7_75t_R n_2275 (.A1(n_2065_o_0),
    .A2(n_2111_o_0),
    .B(n_1928_o_0),
    .Y(n_2275_o_0));
 AOI31xp33_ASAP7_75t_R n_2276 (.A1(n_1936_o_0),
    .A2(n_1932_o_0),
    .A3(net33),
    .B(n_2042_o_0),
    .Y(n_2276_o_0));
 AOI21xp33_ASAP7_75t_R n_2277 (.A1(n_2120_o_0),
    .A2(n_2276_o_0),
    .B(n_1872_o_0),
    .Y(n_2277_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2278 (.A1(net18),
    .A2(n_2275_o_0),
    .B(n_2277_o_0),
    .C(n_2027_o_0),
    .Y(n_2278_o_0));
 OAI21xp33_ASAP7_75t_R n_2279 (.A1(n_2274_o_0),
    .A2(n_1873_o_0),
    .B(n_2278_o_0),
    .Y(n_2279_o_0));
 NAND3xp33_ASAP7_75t_R n_2280 (.A(n_2269_o_0),
    .B(n_1993_o_0),
    .C(n_2279_o_0),
    .Y(n_2280_o_0));
 OAI21xp33_ASAP7_75t_R n_2281 (.A1(n_1993_o_0),
    .A2(n_2262_o_0),
    .B(n_2280_o_0),
    .Y(n_2281_o_0));
 NOR3xp33_ASAP7_75t_R n_2282 (.A(n_1955_o_0),
    .B(n_1932_o_0),
    .C(n_1927_o_0),
    .Y(n_2282_o_0));
 AOI311xp33_ASAP7_75t_R n_2283 (.A1(net33),
    .A2(n_1932_o_0),
    .A3(n_1955_o_0),
    .B(n_2282_o_0),
    .C(n_2186_o_0),
    .Y(n_2283_o_0));
 AOI21xp33_ASAP7_75t_R n_2284 (.A1(n_2067_o_0),
    .A2(n_1998_o_0),
    .B(n_1938_o_0),
    .Y(n_2284_o_0));
 AOI211xp5_ASAP7_75t_R n_2285 (.A1(net8),
    .A2(n_1912_o_0),
    .B(n_2284_o_0),
    .C(net18),
    .Y(n_2285_o_0));
 AOI211xp5_ASAP7_75t_R n_2286 (.A1(n_2283_o_0),
    .A2(net18),
    .B(n_1993_o_0),
    .C(n_2285_o_0),
    .Y(n_2286_o_0));
 OAI22xp33_ASAP7_75t_R n_2287 (.A1(n_2220_o_0),
    .A2(n_2110_o_0),
    .B1(n_2036_o_0),
    .B2(n_1914_o_0),
    .Y(n_2287_o_0));
 OAI211xp5_ASAP7_75t_R n_2288 (.A1(n_2011_o_0),
    .A2(n_1975_o_0),
    .B(n_2182_o_0),
    .C(n_1951_o_0),
    .Y(n_2288_o_0));
 OAI31xp33_ASAP7_75t_R n_2289 (.A1(net98),
    .A2(n_1966_o_0),
    .A3(n_2287_o_0),
    .B(n_2288_o_0),
    .Y(n_2289_o_0));
 NOR2xp33_ASAP7_75t_R n_2290 (.A(net31),
    .B(n_2289_o_0),
    .Y(n_2290_o_0));
 AOI22xp33_ASAP7_75t_R n_2291 (.A1(n_2216_o_0),
    .A2(n_2022_o_0),
    .B1(n_1936_o_0),
    .B2(n_2041_o_0),
    .Y(n_2291_o_0));
 AOI31xp33_ASAP7_75t_R n_2292 (.A1(n_1978_o_0),
    .A2(n_1962_o_0),
    .A3(net33),
    .B(n_1951_o_0),
    .Y(n_2292_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2293 (.A1(n_1975_o_0),
    .A2(n_2011_o_0),
    .B(n_2292_o_0),
    .C(n_1880_o_0),
    .Y(n_2293_o_0));
 INVx1_ASAP7_75t_R n_2294 (.A(n_2293_o_0),
    .Y(n_2294_o_0));
 INVx1_ASAP7_75t_R n_2295 (.A(n_1998_o_0),
    .Y(n_2295_o_0));
 OAI211xp5_ASAP7_75t_R n_2296 (.A1(n_1898_o_0),
    .A2(n_1955_o_0),
    .B(n_2047_o_0),
    .C(n_1938_o_0),
    .Y(n_2296_o_0));
 OAI31xp33_ASAP7_75t_R n_2297 (.A1(n_2164_o_0),
    .A2(n_2295_o_0),
    .A3(net8),
    .B(n_2296_o_0),
    .Y(n_2297_o_0));
 AOI21xp33_ASAP7_75t_R n_2298 (.A1(n_1984_o_0),
    .A2(n_2003_o_0),
    .B(n_1890_o_0),
    .Y(n_2298_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2299 (.A1(n_1973_o_0),
    .A2(net4),
    .B(n_2298_o_0),
    .C(n_1993_o_0),
    .Y(n_2299_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2300 (.A1(n_2297_o_0),
    .A2(net17),
    .B(n_2299_o_0),
    .C(n_1873_o_0),
    .Y(n_2300_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2301 (.A1(net18),
    .A2(n_2291_o_0),
    .B(n_2294_o_0),
    .C(n_2300_o_0),
    .Y(n_2301_o_0));
 OAI31xp33_ASAP7_75t_R n_2302 (.A1(n_2286_o_0),
    .A2(n_2290_o_0),
    .A3(n_1872_o_0),
    .B(n_2301_o_0),
    .Y(n_2302_o_0));
 NAND3xp33_ASAP7_75t_R n_2303 (.A(n_1978_o_0),
    .B(n_2081_o_0),
    .C(net33),
    .Y(n_2303_o_0));
 OAI31xp33_ASAP7_75t_R n_2304 (.A1(net33),
    .A2(n_2295_o_0),
    .A3(n_2170_o_0),
    .B(n_2303_o_0),
    .Y(n_2304_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2305 (.A1(n_2008_o_0),
    .A2(net4),
    .B(n_2220_o_0),
    .C(n_1918_o_0),
    .Y(n_2305_o_0));
 AOI21xp33_ASAP7_75t_R n_2306 (.A1(net18),
    .A2(n_2305_o_0),
    .B(n_1993_o_0),
    .Y(n_2306_o_0));
 OAI21xp33_ASAP7_75t_R n_2307 (.A1(net33),
    .A2(n_2047_o_0),
    .B(n_2182_o_0),
    .Y(n_2307_o_0));
 NAND3xp33_ASAP7_75t_R n_2308 (.A(n_1984_o_0),
    .B(n_1945_o_0),
    .C(n_1938_o_0),
    .Y(n_2308_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2309 (.A1(net4),
    .A2(n_2023_o_0),
    .B(n_2308_o_0),
    .C(n_1890_o_0),
    .Y(n_2309_o_0));
 AOI211xp5_ASAP7_75t_R n_2310 (.A1(n_1890_o_0),
    .A2(n_2307_o_0),
    .B(n_2309_o_0),
    .C(n_1880_o_0),
    .Y(n_2310_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2311 (.A1(net18),
    .A2(n_2304_o_0),
    .B(n_2306_o_0),
    .C(n_2310_o_0),
    .Y(n_2311_o_0));
 AOI21xp33_ASAP7_75t_R n_2312 (.A1(n_1963_o_0),
    .A2(n_2208_o_0),
    .B(n_1890_o_0),
    .Y(n_2312_o_0));
 AOI211xp5_ASAP7_75t_R n_2313 (.A1(n_1890_o_0),
    .A2(n_2139_o_0),
    .B(n_2312_o_0),
    .C(n_1880_o_0),
    .Y(n_2313_o_0));
 NAND2xp33_ASAP7_75t_R n_2314 (.A(n_1941_o_0),
    .B(n_1932_o_0),
    .Y(n_2314_o_0));
 AOI31xp33_ASAP7_75t_R n_2315 (.A1(net4),
    .A2(n_1968_o_0),
    .A3(n_1998_o_0),
    .B(n_1951_o_0),
    .Y(n_2315_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2316 (.A1(n_2314_o_0),
    .A2(n_2075_o_0),
    .B(net8),
    .C(n_2315_o_0),
    .Y(n_2316_o_0));
 OAI31xp33_ASAP7_75t_R n_2317 (.A1(net8),
    .A2(n_2021_o_0),
    .A3(n_1989_o_0),
    .B(n_2063_o_0),
    .Y(n_2317_o_0));
 AOI21xp33_ASAP7_75t_R n_2318 (.A1(n_2316_o_0),
    .A2(n_2317_o_0),
    .B(n_1993_o_0),
    .Y(n_2318_o_0));
 NOR3xp33_ASAP7_75t_R n_2319 (.A(n_2313_o_0),
    .B(n_2318_o_0),
    .C(n_1873_o_0),
    .Y(n_2319_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2320 (.A1(n_2311_o_0),
    .A2(n_1873_o_0),
    .B(n_2319_o_0),
    .C(n_1865_o_0),
    .Y(n_2320_o_0));
 OAI21xp33_ASAP7_75t_R n_2321 (.A1(n_1865_o_0),
    .A2(n_2302_o_0),
    .B(n_2320_o_0),
    .Y(n_2321_o_0));
 NOR2xp33_ASAP7_75t_R n_2322 (.A(n_2200_o_0),
    .B(n_2031_o_0),
    .Y(n_2322_o_0));
 OAI21xp33_ASAP7_75t_R n_2323 (.A1(n_1914_o_0),
    .A2(net4),
    .B(n_1890_o_0),
    .Y(n_2323_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2324 (.A1(n_2119_o_0),
    .A2(n_1955_o_0),
    .B(n_2323_o_0),
    .C(n_1880_o_0),
    .Y(n_2324_o_0));
 AOI31xp33_ASAP7_75t_R n_2325 (.A1(net18),
    .A2(n_2322_o_0),
    .A3(n_2073_o_0),
    .B(n_2324_o_0),
    .Y(n_2325_o_0));
 OAI21xp33_ASAP7_75t_R n_2326 (.A1(n_2072_o_0),
    .A2(n_2021_o_0),
    .B(n_2063_o_0),
    .Y(n_2326_o_0));
 AOI21xp33_ASAP7_75t_R n_2327 (.A1(net8),
    .A2(n_1973_o_0),
    .B(n_2326_o_0),
    .Y(n_2327_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2328 (.A1(n_1898_o_0),
    .A2(n_1936_o_0),
    .B(n_1975_o_0),
    .C(n_1890_o_0),
    .Y(n_2328_o_0));
 AOI21xp33_ASAP7_75t_R n_2329 (.A1(net33),
    .A2(n_1994_o_0),
    .B(n_2328_o_0),
    .Y(n_2329_o_0));
 NOR3xp33_ASAP7_75t_R n_2330 (.A(n_2327_o_0),
    .B(n_2329_o_0),
    .C(net31),
    .Y(n_2330_o_0));
 AOI211xp5_ASAP7_75t_R n_2331 (.A1(n_1932_o_0),
    .A2(n_1937_o_0),
    .B(n_2021_o_0),
    .C(net4),
    .Y(n_2331_o_0));
 AOI211xp5_ASAP7_75t_R n_2332 (.A1(n_1898_o_0),
    .A2(n_1955_o_0),
    .B(n_2049_o_0),
    .C(net33),
    .Y(n_2332_o_0));
 OAI311xp33_ASAP7_75t_R n_2333 (.A1(net33),
    .A2(n_1973_o_0),
    .A3(n_2049_o_0),
    .B1(n_1951_o_0),
    .C1(n_2178_o_0),
    .Y(n_2333_o_0));
 OAI31xp33_ASAP7_75t_R n_2334 (.A1(net17),
    .A2(n_2331_o_0),
    .A3(n_2332_o_0),
    .B(n_2333_o_0),
    .Y(n_2334_o_0));
 INVx1_ASAP7_75t_R n_2335 (.A(n_2284_o_0),
    .Y(n_2335_o_0));
 OAI211xp5_ASAP7_75t_R n_2336 (.A1(net33),
    .A2(n_1942_o_0),
    .B(n_2335_o_0),
    .C(n_1951_o_0),
    .Y(n_2336_o_0));
 NOR3xp33_ASAP7_75t_R n_2337 (.A(n_1951_o_0),
    .B(n_1965_o_0),
    .C(n_2119_o_0),
    .Y(n_2337_o_0));
 NOR3xp33_ASAP7_75t_R n_2338 (.A(n_1951_o_0),
    .B(n_1898_o_0),
    .C(n_1955_o_0),
    .Y(n_2338_o_0));
 OAI22xp33_ASAP7_75t_R n_2339 (.A1(n_2337_o_0),
    .A2(n_2338_o_0),
    .B1(n_1995_o_0),
    .B2(net4),
    .Y(n_2339_o_0));
 NAND3xp33_ASAP7_75t_R n_2340 (.A(n_2336_o_0),
    .B(n_2339_o_0),
    .C(n_1993_o_0),
    .Y(n_2340_o_0));
 OAI211xp5_ASAP7_75t_R n_2341 (.A1(n_1993_o_0),
    .A2(n_2334_o_0),
    .B(n_2340_o_0),
    .C(n_1873_o_0),
    .Y(n_2341_o_0));
 OAI31xp33_ASAP7_75t_R n_2342 (.A1(n_1873_o_0),
    .A2(n_2325_o_0),
    .A3(n_2330_o_0),
    .B(n_2341_o_0),
    .Y(n_2342_o_0));
 NAND2xp33_ASAP7_75t_R n_2343 (.A(n_1962_o_0),
    .B(n_2239_o_0),
    .Y(n_2343_o_0));
 AO21x1_ASAP7_75t_R n_2344 (.A1(n_1955_o_0),
    .A2(n_1898_o_0),
    .B(n_2132_o_0),
    .Y(n_2344_o_0));
 OAI21xp33_ASAP7_75t_R n_2345 (.A1(n_1986_o_0),
    .A2(n_2181_o_0),
    .B(n_1993_o_0),
    .Y(n_2345_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2346 (.A1(n_1932_o_0),
    .A2(n_1914_o_0),
    .B(n_2153_o_0),
    .C(n_2345_o_0),
    .Y(n_2346_o_0));
 AOI31xp33_ASAP7_75t_R n_2347 (.A1(n_2343_o_0),
    .A2(n_2344_o_0),
    .A3(net31),
    .B(n_2346_o_0),
    .Y(n_2347_o_0));
 NAND2xp33_ASAP7_75t_R n_2348 (.A(n_2220_o_0),
    .B(n_2208_o_0),
    .Y(n_2348_o_0));
 OAI211xp5_ASAP7_75t_R n_2349 (.A1(n_2220_o_0),
    .A2(n_2110_o_0),
    .B(n_2105_o_0),
    .C(n_1993_o_0),
    .Y(n_2349_o_0));
 OAI21xp33_ASAP7_75t_R n_2350 (.A1(n_1993_o_0),
    .A2(n_2348_o_0),
    .B(n_2349_o_0),
    .Y(n_2350_o_0));
 OAI21xp33_ASAP7_75t_R n_2351 (.A1(net18),
    .A2(n_2350_o_0),
    .B(n_1873_o_0),
    .Y(n_2351_o_0));
 OAI31xp33_ASAP7_75t_R n_2352 (.A1(net33),
    .A2(n_2021_o_0),
    .A3(n_2049_o_0),
    .B(n_2215_o_0),
    .Y(n_2352_o_0));
 NAND3xp33_ASAP7_75t_R n_2353 (.A(n_1995_o_0),
    .B(n_2009_o_0),
    .C(n_1927_o_0),
    .Y(n_2353_o_0));
 OAI211xp5_ASAP7_75t_R n_2354 (.A1(net33),
    .A2(n_1917_o_0),
    .B(n_2353_o_0),
    .C(net31),
    .Y(n_2354_o_0));
 OAI211xp5_ASAP7_75t_R n_2355 (.A1(n_1880_o_0),
    .A2(n_2352_o_0),
    .B(n_2354_o_0),
    .C(net17),
    .Y(n_2355_o_0));
 OAI211xp5_ASAP7_75t_R n_2356 (.A1(n_1898_o_0),
    .A2(n_1915_o_0),
    .B(n_1998_o_0),
    .C(n_1938_o_0),
    .Y(n_2356_o_0));
 OAI31xp33_ASAP7_75t_R n_2357 (.A1(n_2008_o_0),
    .A2(n_1973_o_0),
    .A3(net4),
    .B(n_2356_o_0),
    .Y(n_2357_o_0));
 INVx1_ASAP7_75t_R n_2358 (.A(n_2240_o_0),
    .Y(n_2358_o_0));
 NOR3xp33_ASAP7_75t_R n_2359 (.A(n_2168_o_0),
    .B(n_1880_o_0),
    .C(n_2358_o_0),
    .Y(n_2359_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2360 (.A1(n_1880_o_0),
    .A2(n_2357_o_0),
    .B(n_2359_o_0),
    .C(n_1890_o_0),
    .Y(n_2360_o_0));
 AOI31xp33_ASAP7_75t_R n_2361 (.A1(n_1872_o_0),
    .A2(n_2355_o_0),
    .A3(n_2360_o_0),
    .B(n_2027_o_0),
    .Y(n_2361_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2362 (.A1(net18),
    .A2(n_2347_o_0),
    .B(n_2351_o_0),
    .C(n_2361_o_0),
    .Y(n_2362_o_0));
 OAI21xp33_ASAP7_75t_R n_2363 (.A1(n_1865_o_0),
    .A2(n_2342_o_0),
    .B(n_2362_o_0),
    .Y(n_2363_o_0));
 XOR2xp5_ASAP7_75t_R n_2364 (.A(_00453_),
    .B(_00995_),
    .Y(n_2364_o_0));
 XOR2xp5_ASAP7_75t_R n_2365 (.A(_00891_),
    .B(n_2364_o_0),
    .Y(n_2365_o_0));
 XNOR2xp5_ASAP7_75t_R n_2366 (.A(_00923_),
    .B(n_2365_o_0),
    .Y(n_2366_o_0));
 INVx1_ASAP7_75t_R n_2367 (.A(n_2366_o_0),
    .Y(n_2367_o_0));
 XNOR2xp5_ASAP7_75t_R n_2368 (.A(_00955_),
    .B(n_2367_o_0),
    .Y(n_2368_o_0));
 INVx1_ASAP7_75t_R n_2369 (.A(_00987_),
    .Y(n_2369_o_0));
 NOR2xp33_ASAP7_75t_R n_2370 (.A(n_2369_o_0),
    .B(n_2368_o_0),
    .Y(n_2370_o_0));
 NOR2xp33_ASAP7_75t_R n_2371 (.A(key[31]),
    .B(n_827_o_0),
    .Y(n_2371_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2372 (.A1(n_2368_o_0),
    .A2(n_2369_o_0),
    .B(n_2370_o_0),
    .C(n_827_o_0),
    .D(n_2371_o_0),
    .Y(n_2372_o_0));
 INVx1_ASAP7_75t_R n_2373 (.A(n_2372_o_0),
    .Y(n_2373_o_0));
 INVx1_ASAP7_75t_R n_2374 (.A(_00986_),
    .Y(n_2374_o_0));
 XOR2xp5_ASAP7_75t_R n_2375 (.A(_00452_),
    .B(_00994_),
    .Y(n_2375_o_0));
 XNOR2xp5_ASAP7_75t_R n_2376 (.A(_00890_),
    .B(n_2375_o_0),
    .Y(n_2376_o_0));
 XNOR2xp5_ASAP7_75t_R n_2377 (.A(_00922_),
    .B(n_2376_o_0),
    .Y(n_2377_o_0));
 INVx1_ASAP7_75t_R n_2378 (.A(_00954_),
    .Y(n_2378_o_0));
 NAND2xp33_ASAP7_75t_R n_2379 (.A(n_2378_o_0),
    .B(n_2377_o_0),
    .Y(n_2379_o_0));
 OAI21xp33_ASAP7_75t_R n_2380 (.A1(n_2377_o_0),
    .A2(n_2378_o_0),
    .B(n_2379_o_0),
    .Y(n_2380_o_0));
 INVx1_ASAP7_75t_R n_2381 (.A(n_2380_o_0),
    .Y(n_2381_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2382 (.A1(n_2378_o_0),
    .A2(n_2377_o_0),
    .B(n_2379_o_0),
    .C(n_2374_o_0),
    .Y(n_2382_o_0));
 NOR2xp33_ASAP7_75t_R n_2383 (.A(key[30]),
    .B(n_827_o_0),
    .Y(n_2383_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2384 (.A1(n_2374_o_0),
    .A2(n_2381_o_0),
    .B(n_2382_o_0),
    .C(n_827_o_0),
    .D(n_2383_o_0),
    .Y(n_2384_o_0));
 INVx1_ASAP7_75t_R n_2385 (.A(n_2384_o_0),
    .Y(n_2385_o_0));
 INVx1_ASAP7_75t_R n_2386 (.A(_00953_),
    .Y(n_2386_o_0));
 XOR2xp5_ASAP7_75t_R n_2387 (.A(_00451_),
    .B(_00993_),
    .Y(n_2387_o_0));
 XNOR2xp5_ASAP7_75t_R n_2388 (.A(_00889_),
    .B(n_2387_o_0),
    .Y(n_2388_o_0));
 XNOR2xp5_ASAP7_75t_R n_2389 (.A(_00921_),
    .B(n_2388_o_0),
    .Y(n_2389_o_0));
 NOR2xp33_ASAP7_75t_R n_2390 (.A(n_2386_o_0),
    .B(n_2389_o_0),
    .Y(n_2390_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2391 (.A1(n_2386_o_0),
    .A2(n_2389_o_0),
    .B(n_2390_o_0),
    .C(_00985_),
    .Y(n_2391_o_0));
 NAND2xp33_ASAP7_75t_R n_2392 (.A(n_2386_o_0),
    .B(n_2389_o_0),
    .Y(n_2392_o_0));
 INVx1_ASAP7_75t_R n_2393 (.A(_00985_),
    .Y(n_2393_o_0));
 OAI211xp5_ASAP7_75t_R n_2394 (.A1(n_2386_o_0),
    .A2(n_2389_o_0),
    .B(n_2392_o_0),
    .C(n_2393_o_0),
    .Y(n_2394_o_0));
 AND2x2_ASAP7_75t_R n_2395 (.A(key[29]),
    .B(ld),
    .Y(n_2395_o_0));
 AOI31xp33_ASAP7_75t_R n_2396 (.A1(n_827_o_0),
    .A2(n_2391_o_0),
    .A3(n_2394_o_0),
    .B(n_2395_o_0),
    .Y(n_2396_o_0));
 NOR2xp33_ASAP7_75t_R n_2397 (.A(_00449_),
    .B(_00991_),
    .Y(n_2397_o_0));
 AND2x2_ASAP7_75t_R n_2398 (.A(_00449_),
    .B(_00991_),
    .Y(n_2398_o_0));
 INVx1_ASAP7_75t_R n_2399 (.A(_00919_),
    .Y(n_2399_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2400 (.A1(_00449_),
    .A2(_00991_),
    .B(n_2397_o_0),
    .C(_00887_),
    .Y(n_2400_o_0));
 OAI311xp33_ASAP7_75t_R n_2401 (.A1(_00887_),
    .A2(n_2397_o_0),
    .A3(n_2398_o_0),
    .B1(n_2399_o_0),
    .C1(n_2400_o_0),
    .Y(n_2401_o_0));
 INVx1_ASAP7_75t_R n_2402 (.A(_00887_),
    .Y(n_2402_o_0));
 XOR2xp5_ASAP7_75t_R n_2403 (.A(_00449_),
    .B(_00991_),
    .Y(n_2403_o_0));
 INVx1_ASAP7_75t_R n_2404 (.A(n_2400_o_0),
    .Y(n_2404_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2405 (.A1(n_2402_o_0),
    .A2(n_2403_o_0),
    .B(n_2404_o_0),
    .C(_00919_),
    .Y(n_2405_o_0));
 INVx1_ASAP7_75t_R n_2406 (.A(_00951_),
    .Y(n_2406_o_0));
 NAND2xp33_ASAP7_75t_R n_2407 (.A(n_2402_o_0),
    .B(n_2403_o_0),
    .Y(n_2407_o_0));
 OAI21xp33_ASAP7_75t_R n_2408 (.A1(n_2403_o_0),
    .A2(n_2402_o_0),
    .B(n_2407_o_0),
    .Y(n_2408_o_0));
 OAI211xp5_ASAP7_75t_R n_2409 (.A1(n_2408_o_0),
    .A2(_00919_),
    .B(n_2405_o_0),
    .C(n_2406_o_0),
    .Y(n_2409_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2410 (.A1(n_2401_o_0),
    .A2(n_2405_o_0),
    .B(n_2406_o_0),
    .C(n_2409_o_0),
    .D(_00983_),
    .Y(n_2410_o_0));
 INVx1_ASAP7_75t_R n_2411 (.A(_00983_),
    .Y(n_2411_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2412 (.A1(n_2400_o_0),
    .A2(n_2407_o_0),
    .B(n_2399_o_0),
    .C(n_2401_o_0),
    .D(n_2406_o_0),
    .Y(n_2412_o_0));
 AOI311xp33_ASAP7_75t_R n_2413 (.A1(n_2406_o_0),
    .A2(n_2401_o_0),
    .A3(n_2405_o_0),
    .B(n_2411_o_0),
    .C(n_2412_o_0),
    .Y(n_2413_o_0));
 OR2x2_ASAP7_75t_R n_2414 (.A(key[27]),
    .B(n_827_o_0),
    .Y(n_2414_o_0));
 OAI31xp67_ASAP7_75t_R n_2415 (.A1(ld),
    .A2(n_2410_o_0),
    .A3(n_2413_o_0),
    .B(n_2414_o_0),
    .Y(n_2415_o_0));
 NAND2xp33_ASAP7_75t_R n_2416 (.A(_00446_),
    .B(_00988_),
    .Y(n_2416_o_0));
 INVx1_ASAP7_75t_R n_2417 (.A(_00884_),
    .Y(n_2417_o_0));
 OAI211xp5_ASAP7_75t_R n_2418 (.A1(_00446_),
    .A2(_00988_),
    .B(n_2416_o_0),
    .C(n_2417_o_0),
    .Y(n_2418_o_0));
 NOR2xp33_ASAP7_75t_R n_2419 (.A(_00446_),
    .B(_00988_),
    .Y(n_2419_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2420 (.A1(_00446_),
    .A2(_00988_),
    .B(n_2419_o_0),
    .C(_00884_),
    .Y(n_2420_o_0));
 INVx1_ASAP7_75t_R n_2421 (.A(_00916_),
    .Y(n_2421_o_0));
 AOI21xp33_ASAP7_75t_R n_2422 (.A1(n_2418_o_0),
    .A2(n_2420_o_0),
    .B(n_2421_o_0),
    .Y(n_2422_o_0));
 AOI21xp33_ASAP7_75t_R n_2423 (.A1(_00446_),
    .A2(_00988_),
    .B(n_2419_o_0),
    .Y(n_2423_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2424 (.A1(_00446_),
    .A2(_00988_),
    .B(n_2416_o_0),
    .C(n_2417_o_0),
    .Y(n_2424_o_0));
 AOI211xp5_ASAP7_75t_R n_2425 (.A1(n_2423_o_0),
    .A2(n_2417_o_0),
    .B(_00916_),
    .C(n_2424_o_0),
    .Y(n_2425_o_0));
 OAI21xp33_ASAP7_75t_R n_2426 (.A1(n_2422_o_0),
    .A2(n_2425_o_0),
    .B(_00948_),
    .Y(n_2426_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2427 (.A1(n_2423_o_0),
    .A2(n_2417_o_0),
    .B(n_2424_o_0),
    .C(_00916_),
    .Y(n_2427_o_0));
 INVx1_ASAP7_75t_R n_2428 (.A(n_2416_o_0),
    .Y(n_2428_o_0));
 OAI311xp33_ASAP7_75t_R n_2429 (.A1(_00884_),
    .A2(n_2428_o_0),
    .A3(n_2419_o_0),
    .B1(n_2421_o_0),
    .C1(n_2420_o_0),
    .Y(n_2429_o_0));
 INVx1_ASAP7_75t_R n_2430 (.A(_00948_),
    .Y(n_2430_o_0));
 NAND3xp33_ASAP7_75t_R n_2431 (.A(n_2427_o_0),
    .B(n_2429_o_0),
    .C(n_2430_o_0),
    .Y(n_2431_o_0));
 INVx1_ASAP7_75t_R n_2432 (.A(_00980_),
    .Y(n_2432_o_0));
 AOI21xp33_ASAP7_75t_R n_2433 (.A1(n_2426_o_0),
    .A2(n_2431_o_0),
    .B(n_2432_o_0),
    .Y(n_2433_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2434 (.A1(n_2418_o_0),
    .A2(n_2420_o_0),
    .B(n_2421_o_0),
    .C(n_2429_o_0),
    .D(n_2430_o_0),
    .Y(n_2434_o_0));
 AOI311xp33_ASAP7_75t_R n_2435 (.A1(n_2430_o_0),
    .A2(n_2429_o_0),
    .A3(n_2427_o_0),
    .B(_00980_),
    .C(n_2434_o_0),
    .Y(n_2435_o_0));
 NAND2xp33_ASAP7_75t_R n_2436 (.A(key[24]),
    .B(ld),
    .Y(n_2436_o_0));
 OAI31xp67_ASAP7_75t_R n_2437 (.A1(n_2435_o_0),
    .A2(n_2433_o_0),
    .A3(ld),
    .B(n_2436_o_0),
    .Y(n_2437_o_0));
 INVx1_ASAP7_75t_R n_2438 (.A(_00885_),
    .Y(n_2438_o_0));
 NOR2xp33_ASAP7_75t_R n_2439 (.A(_00447_),
    .B(_00989_),
    .Y(n_2439_o_0));
 AOI21xp33_ASAP7_75t_R n_2440 (.A1(_00447_),
    .A2(_00989_),
    .B(n_2439_o_0),
    .Y(n_2440_o_0));
 NAND2xp33_ASAP7_75t_R n_2441 (.A(_00447_),
    .B(_00989_),
    .Y(n_2441_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2442 (.A1(_00447_),
    .A2(_00989_),
    .B(n_2441_o_0),
    .C(n_2438_o_0),
    .Y(n_2442_o_0));
 AOI211xp5_ASAP7_75t_R n_2443 (.A1(n_2440_o_0),
    .A2(n_2438_o_0),
    .B(_00917_),
    .C(n_2442_o_0),
    .Y(n_2443_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2444 (.A1(n_2438_o_0),
    .A2(n_2440_o_0),
    .B(n_2442_o_0),
    .C(_00917_),
    .D(n_2443_o_0),
    .Y(n_2444_o_0));
 INVx1_ASAP7_75t_R n_2445 (.A(_00949_),
    .Y(n_2445_o_0));
 INVx1_ASAP7_75t_R n_2446 (.A(n_2441_o_0),
    .Y(n_2446_o_0));
 INVx1_ASAP7_75t_R n_2447 (.A(_00917_),
    .Y(n_2447_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2448 (.A1(_00447_),
    .A2(_00989_),
    .B(n_2439_o_0),
    .C(_00885_),
    .Y(n_2448_o_0));
 OAI311xp33_ASAP7_75t_R n_2449 (.A1(_00885_),
    .A2(n_2446_o_0),
    .A3(n_2439_o_0),
    .B1(n_2447_o_0),
    .C1(n_2448_o_0),
    .Y(n_2449_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2450 (.A1(n_2440_o_0),
    .A2(n_2438_o_0),
    .B(n_2442_o_0),
    .C(_00917_),
    .Y(n_2450_o_0));
 AOI21xp33_ASAP7_75t_R n_2451 (.A1(n_2449_o_0),
    .A2(n_2450_o_0),
    .B(n_2445_o_0),
    .Y(n_2451_o_0));
 AOI211xp5_ASAP7_75t_R n_2452 (.A1(n_2444_o_0),
    .A2(n_2445_o_0),
    .B(_00981_),
    .C(n_2451_o_0),
    .Y(n_2452_o_0));
 OAI211xp5_ASAP7_75t_R n_2453 (.A1(_00447_),
    .A2(_00989_),
    .B(n_2441_o_0),
    .C(n_2438_o_0),
    .Y(n_2453_o_0));
 OAI21xp33_ASAP7_75t_R n_2454 (.A1(n_2438_o_0),
    .A2(n_2440_o_0),
    .B(n_2453_o_0),
    .Y(n_2454_o_0));
 OAI211xp5_ASAP7_75t_R n_2455 (.A1(n_2454_o_0),
    .A2(_00917_),
    .B(n_2450_o_0),
    .C(n_2445_o_0),
    .Y(n_2455_o_0));
 INVx1_ASAP7_75t_R n_2456 (.A(_00981_),
    .Y(n_2456_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2457 (.A1(n_2449_o_0),
    .A2(n_2450_o_0),
    .B(n_2445_o_0),
    .C(n_2455_o_0),
    .D(n_2456_o_0),
    .Y(n_2457_o_0));
 NAND2xp33_ASAP7_75t_R n_2458 (.A(key[25]),
    .B(ld),
    .Y(n_2458_o_0));
 OAI31xp67_ASAP7_75t_R n_2459 (.A1(n_2452_o_0),
    .A2(ld),
    .A3(n_2457_o_0),
    .B(n_2458_o_0),
    .Y(n_2459_o_0));
 NAND2xp33_ASAP7_75t_R n_2460 (.A(n_2437_o_0),
    .B(n_2459_o_0),
    .Y(n_2460_o_0));
 INVx1_ASAP7_75t_R n_2461 (.A(n_2460_o_0),
    .Y(n_2461_o_0));
 INVx1_ASAP7_75t_R n_2462 (.A(_00950_),
    .Y(n_2462_o_0));
 INVx1_ASAP7_75t_R n_2463 (.A(_00918_),
    .Y(n_2463_o_0));
 INVx1_ASAP7_75t_R n_2464 (.A(_00886_),
    .Y(n_2464_o_0));
 XNOR2xp5_ASAP7_75t_R n_2465 (.A(_00448_),
    .B(_00990_),
    .Y(n_2465_o_0));
 XNOR2xp5_ASAP7_75t_R n_2466 (.A(n_2464_o_0),
    .B(n_2465_o_0),
    .Y(n_2466_o_0));
 INVx1_ASAP7_75t_R n_2467 (.A(_00990_),
    .Y(n_2467_o_0));
 NAND2xp33_ASAP7_75t_R n_2468 (.A(_00448_),
    .B(n_2467_o_0),
    .Y(n_2468_o_0));
 OAI211xp5_ASAP7_75t_R n_2469 (.A1(_00448_),
    .A2(n_2467_o_0),
    .B(n_2468_o_0),
    .C(_00886_),
    .Y(n_2469_o_0));
 NOR2xp33_ASAP7_75t_R n_2470 (.A(_00448_),
    .B(n_2467_o_0),
    .Y(n_2470_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2471 (.A1(_00448_),
    .A2(n_2467_o_0),
    .B(n_2470_o_0),
    .C(n_2464_o_0),
    .Y(n_2471_o_0));
 AOI21xp33_ASAP7_75t_R n_2472 (.A1(n_2469_o_0),
    .A2(n_2471_o_0),
    .B(n_2463_o_0),
    .Y(n_2472_o_0));
 AOI21xp33_ASAP7_75t_R n_2473 (.A1(n_2463_o_0),
    .A2(n_2466_o_0),
    .B(n_2472_o_0),
    .Y(n_2473_o_0));
 OAI211xp5_ASAP7_75t_R n_2474 (.A1(_00886_),
    .A2(n_2465_o_0),
    .B(n_2469_o_0),
    .C(n_2463_o_0),
    .Y(n_2474_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2475 (.A1(n_2469_o_0),
    .A2(n_2471_o_0),
    .B(n_2463_o_0),
    .C(n_2474_o_0),
    .D(n_2462_o_0),
    .Y(n_2475_o_0));
 AOI21xp33_ASAP7_75t_R n_2476 (.A1(n_2462_o_0),
    .A2(n_2473_o_0),
    .B(n_2475_o_0),
    .Y(n_2476_o_0));
 NOR2xp33_ASAP7_75t_R n_2477 (.A(_00886_),
    .B(n_2465_o_0),
    .Y(n_2477_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2478 (.A1(_00886_),
    .A2(n_2465_o_0),
    .B(n_2477_o_0),
    .C(_00918_),
    .Y(n_2478_o_0));
 INVx1_ASAP7_75t_R n_2479 (.A(n_2469_o_0),
    .Y(n_2479_o_0));
 OAI311xp33_ASAP7_75t_R n_2480 (.A1(_00918_),
    .A2(n_2479_o_0),
    .A3(n_2477_o_0),
    .B1(n_2462_o_0),
    .C1(n_2478_o_0),
    .Y(n_2480_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2481 (.A1(n_2474_o_0),
    .A2(n_2478_o_0),
    .B(n_2462_o_0),
    .C(n_2480_o_0),
    .D(_00982_),
    .Y(n_2481_o_0));
 NAND2xp33_ASAP7_75t_R n_2482 (.A(key[26]),
    .B(ld),
    .Y(n_2482_o_0));
 INVx1_ASAP7_75t_R n_2483 (.A(n_2482_o_0),
    .Y(n_2483_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2484 (.A1(_00982_),
    .A2(n_2476_o_0),
    .B(n_2481_o_0),
    .C(n_827_o_0),
    .D(n_2483_o_0),
    .Y(n_2484_o_0));
 NAND2xp33_ASAP7_75t_R n_2485 (.A(n_2415_o_0),
    .B(n_2484_o_0),
    .Y(n_2485_o_0));
 OAI32xp33_ASAP7_75t_R n_2486 (.A1(net52),
    .A2(n_2461_o_0),
    .A3(net21),
    .B1(n_2485_o_0),
    .B2(net100),
    .Y(n_2486_o_0));
 INVx1_ASAP7_75t_R n_2487 (.A(_00982_),
    .Y(n_2487_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2488 (.A1(n_2473_o_0),
    .A2(n_2462_o_0),
    .B(n_2475_o_0),
    .C(n_2487_o_0),
    .Y(n_2488_o_0));
 AOI211xp5_ASAP7_75t_R n_2489 (.A1(_00886_),
    .A2(n_2465_o_0),
    .B(n_2477_o_0),
    .C(_00918_),
    .Y(n_2489_o_0));
 OAI21xp33_ASAP7_75t_R n_2490 (.A1(n_2472_o_0),
    .A2(n_2489_o_0),
    .B(_00950_),
    .Y(n_2490_o_0));
 OAI311xp33_ASAP7_75t_R n_2491 (.A1(_00950_),
    .A2(n_2489_o_0),
    .A3(n_2472_o_0),
    .B1(_00982_),
    .C1(n_2490_o_0),
    .Y(n_2491_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2492 (.A1(n_2491_o_0),
    .A2(n_2488_o_0),
    .B(ld),
    .C(n_2482_o_0),
    .Y(n_2492_o_0));
 NAND2xp33_ASAP7_75t_R n_2493 (.A(n_2418_o_0),
    .B(n_2420_o_0),
    .Y(n_2493_o_0));
 AOI211xp5_ASAP7_75t_R n_2494 (.A1(n_2493_o_0),
    .A2(_00916_),
    .B(_00948_),
    .C(n_2425_o_0),
    .Y(n_2494_o_0));
 OAI21xp33_ASAP7_75t_R n_2495 (.A1(n_2434_o_0),
    .A2(n_2494_o_0),
    .B(_00980_),
    .Y(n_2495_o_0));
 OAI311xp33_ASAP7_75t_R n_2496 (.A1(_00948_),
    .A2(n_2425_o_0),
    .A3(n_2422_o_0),
    .B1(n_2432_o_0),
    .C1(n_2426_o_0),
    .Y(n_2496_o_0));
 INVx1_ASAP7_75t_R n_2497 (.A(n_2436_o_0),
    .Y(n_2497_o_0));
 AOI31xp67_ASAP7_75t_R n_2498 (.A1(n_827_o_0),
    .A2(n_2495_o_0),
    .A3(n_2496_o_0),
    .B(n_2497_o_0),
    .Y(n_2498_o_0));
 NOR3xp33_ASAP7_75t_R n_2499 (.A(n_2492_o_0),
    .B(n_2415_o_0),
    .C(n_2498_o_0),
    .Y(n_2499_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2500 (.A1(n_2444_o_0),
    .A2(n_2445_o_0),
    .B(n_2451_o_0),
    .C(_00981_),
    .Y(n_2500_o_0));
 AOI21xp33_ASAP7_75t_R n_2501 (.A1(n_2453_o_0),
    .A2(n_2448_o_0),
    .B(n_2447_o_0),
    .Y(n_2501_o_0));
 OAI21xp33_ASAP7_75t_R n_2502 (.A1(n_2501_o_0),
    .A2(n_2443_o_0),
    .B(_00949_),
    .Y(n_2502_o_0));
 OAI311xp33_ASAP7_75t_R n_2503 (.A1(_00949_),
    .A2(n_2443_o_0),
    .A3(n_2501_o_0),
    .B1(n_2456_o_0),
    .C1(n_2502_o_0),
    .Y(n_2503_o_0));
 INVx1_ASAP7_75t_R n_2504 (.A(n_2458_o_0),
    .Y(n_2504_o_0));
 AOI31xp33_ASAP7_75t_R n_2505 (.A1(n_827_o_0),
    .A2(n_2500_o_0),
    .A3(n_2503_o_0),
    .B(n_2504_o_0),
    .Y(n_2505_o_0));
 NAND2xp33_ASAP7_75t_R n_2506 (.A(n_2498_o_0),
    .B(n_2505_o_0),
    .Y(n_2506_o_0));
 OA31x2_ASAP7_75t_R n_2507 (.A1(ld),
    .A2(n_2410_o_0),
    .A3(n_2413_o_0),
    .B1(n_2414_o_0),
    .Y(n_2507_o_0));
 NOR3xp33_ASAP7_75t_R n_2508 (.A(n_2506_o_0),
    .B(n_2507_o_0),
    .C(net75),
    .Y(n_2508_o_0));
 NOR3xp33_ASAP7_75t_R n_2509 (.A(n_2486_o_0),
    .B(n_2499_o_0),
    .C(n_2508_o_0),
    .Y(n_2509_o_0));
 NAND2xp5_ASAP7_75t_R n_2510 (.A(n_2498_o_0),
    .B(n_2459_o_0),
    .Y(n_2510_o_0));
 INVx1_ASAP7_75t_R n_2511 (.A(n_2510_o_0),
    .Y(n_2511_o_0));
 OAI21xp33_ASAP7_75t_R n_2512 (.A1(n_2484_o_0),
    .A2(n_2511_o_0),
    .B(n_2507_o_0),
    .Y(n_2512_o_0));
 AOI21xp33_ASAP7_75t_R n_2513 (.A1(net21),
    .A2(n_2511_o_0),
    .B(n_2512_o_0),
    .Y(n_2513_o_0));
 AOI21xp33_ASAP7_75t_R n_2514 (.A1(n_2498_o_0),
    .A2(net21),
    .B(n_2507_o_0),
    .Y(n_2514_o_0));
 NOR3xp33_ASAP7_75t_R n_2515 (.A(n_2513_o_0),
    .B(n_2396_o_0),
    .C(n_2514_o_0),
    .Y(n_2515_o_0));
 XNOR2xp5_ASAP7_75t_R n_2516 (.A(_00450_),
    .B(_00992_),
    .Y(n_2516_o_0));
 XNOR2xp5_ASAP7_75t_R n_2517 (.A(_00888_),
    .B(n_2516_o_0),
    .Y(n_2517_o_0));
 NAND2xp33_ASAP7_75t_R n_2518 (.A(_00920_),
    .B(n_2517_o_0),
    .Y(n_2518_o_0));
 OA21x2_ASAP7_75t_R n_2519 (.A1(_00920_),
    .A2(n_2517_o_0),
    .B(n_2518_o_0),
    .Y(n_2519_o_0));
 INVx1_ASAP7_75t_R n_2520 (.A(_00952_),
    .Y(n_2520_o_0));
 INVx1_ASAP7_75t_R n_2521 (.A(_00984_),
    .Y(n_2521_o_0));
 OAI211xp5_ASAP7_75t_R n_2522 (.A1(n_2517_o_0),
    .A2(_00920_),
    .B(n_2518_o_0),
    .C(n_2520_o_0),
    .Y(n_2522_o_0));
 OAI211xp5_ASAP7_75t_R n_2523 (.A1(n_2519_o_0),
    .A2(n_2520_o_0),
    .B(n_2521_o_0),
    .C(n_2522_o_0),
    .Y(n_2523_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2524 (.A1(n_2517_o_0),
    .A2(_00920_),
    .B(n_2518_o_0),
    .C(n_2520_o_0),
    .Y(n_2524_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2525 (.A1(n_2519_o_0),
    .A2(n_2520_o_0),
    .B(n_2524_o_0),
    .C(_00984_),
    .Y(n_2525_o_0));
 AND2x2_ASAP7_75t_R n_2526 (.A(key[28]),
    .B(ld),
    .Y(n_2526_o_0));
 AO31x2_ASAP7_75t_R n_2527 (.A1(n_2523_o_0),
    .A2(n_2525_o_0),
    .A3(n_827_o_0),
    .B(n_2526_o_0),
    .Y(n_2527_o_0));
 AOI211xp5_ASAP7_75t_R n_2528 (.A1(n_2396_o_0),
    .A2(n_2509_o_0),
    .B(n_2515_o_0),
    .C(n_2527_o_0),
    .Y(n_2528_o_0));
 AOI21xp33_ASAP7_75t_R n_2529 (.A1(n_2386_o_0),
    .A2(n_2389_o_0),
    .B(n_2390_o_0),
    .Y(n_2529_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2530 (.A1(n_2386_o_0),
    .A2(n_2389_o_0),
    .B(n_2392_o_0),
    .C(n_2393_o_0),
    .Y(n_2530_o_0));
 NOR2xp33_ASAP7_75t_R n_2531 (.A(key[29]),
    .B(n_827_o_0),
    .Y(n_2531_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2532 (.A1(n_2393_o_0),
    .A2(n_2529_o_0),
    .B(n_2530_o_0),
    .C(n_827_o_0),
    .D(n_2531_o_0),
    .Y(n_2532_o_0));
 XNOR2xp5_ASAP7_75t_R n_2533 (.A(_00982_),
    .B(n_2476_o_0),
    .Y(n_2533_o_0));
 INVx1_ASAP7_75t_R n_2534 (.A(key[25]),
    .Y(n_2534_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2535 (.A1(n_2455_o_0),
    .A2(n_2502_o_0),
    .B(n_2456_o_0),
    .C(n_2503_o_0),
    .Y(n_2535_o_0));
 AOI21xp33_ASAP7_75t_R n_2536 (.A1(n_2445_o_0),
    .A2(n_2444_o_0),
    .B(n_2451_o_0),
    .Y(n_2536_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2537 (.A1(n_2536_o_0),
    .A2(n_2456_o_0),
    .B(n_2457_o_0),
    .C(n_2504_o_0),
    .Y(n_2537_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2538 (.A1(n_2534_o_0),
    .A2(ld),
    .B(n_2535_o_0),
    .C(n_2537_o_0),
    .D(n_2498_o_0),
    .Y(n_2538_o_0));
 AOI21xp33_ASAP7_75t_R n_2539 (.A1(n_2456_o_0),
    .A2(n_2536_o_0),
    .B(n_2457_o_0),
    .Y(n_2539_o_0));
 AOI211xp5_ASAP7_75t_R n_2540 (.A1(n_2539_o_0),
    .A2(n_827_o_0),
    .B(n_2437_o_0),
    .C(n_2504_o_0),
    .Y(n_2540_o_0));
 NOR2xp33_ASAP7_75t_R n_2541 (.A(key[26]),
    .B(n_827_o_0),
    .Y(n_2541_o_0));
 INVx1_ASAP7_75t_R n_2542 (.A(n_2541_o_0),
    .Y(n_2542_o_0));
 OAI221xp5_ASAP7_75t_R n_2543 (.A1(ld),
    .A2(n_2533_o_0),
    .B1(n_2538_o_0),
    .B2(n_2540_o_0),
    .C(n_2542_o_0),
    .Y(n_2543_o_0));
 AND2x2_ASAP7_75t_R n_2544 (.A(n_2543_o_0),
    .B(n_2507_o_0),
    .Y(n_2544_o_0));
 NAND2xp33_ASAP7_75t_R n_2545 (.A(n_2484_o_0),
    .B(n_2460_o_0),
    .Y(n_2545_o_0));
 OAI21xp33_ASAP7_75t_R n_2546 (.A1(_00982_),
    .A2(n_2476_o_0),
    .B(n_2491_o_0),
    .Y(n_2546_o_0));
 NAND3xp33_ASAP7_75t_R n_2547 (.A(n_2459_o_0),
    .B(n_2498_o_0),
    .C(n_2482_o_0),
    .Y(n_2547_o_0));
 AO21x1_ASAP7_75t_R n_2548 (.A1(n_827_o_0),
    .A2(n_2546_o_0),
    .B(n_2547_o_0),
    .Y(n_2548_o_0));
 OAI211xp5_ASAP7_75t_R n_2549 (.A1(net102),
    .A2(net21),
    .B(n_2548_o_0),
    .C(n_2415_o_0),
    .Y(n_2549_o_0));
 INVx1_ASAP7_75t_R n_2550 (.A(n_2549_o_0),
    .Y(n_2550_o_0));
 AOI21xp33_ASAP7_75t_R n_2551 (.A1(n_2544_o_0),
    .A2(n_2545_o_0),
    .B(n_2550_o_0),
    .Y(n_2551_o_0));
 NAND2xp33_ASAP7_75t_R n_2552 (.A(n_2498_o_0),
    .B(net75),
    .Y(n_2552_o_0));
 AOI21xp33_ASAP7_75t_R n_2553 (.A1(net101),
    .A2(n_2460_o_0),
    .B(n_2415_o_0),
    .Y(n_2553_o_0));
 OAI21xp33_ASAP7_75t_R n_2554 (.A1(n_2459_o_0),
    .A2(n_2484_o_0),
    .B(n_2415_o_0),
    .Y(n_2554_o_0));
 AOI21xp33_ASAP7_75t_R n_2555 (.A1(n_827_o_0),
    .A2(n_2546_o_0),
    .B(n_2547_o_0),
    .Y(n_2555_o_0));
 OAI21xp33_ASAP7_75t_R n_2556 (.A1(n_2554_o_0),
    .A2(n_2555_o_0),
    .B(n_2396_o_0),
    .Y(n_2556_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2557 (.A1(n_2552_o_0),
    .A2(n_2553_o_0),
    .B(n_2556_o_0),
    .C(n_2527_o_0),
    .Y(n_2557_o_0));
 AOI21xp33_ASAP7_75t_R n_2558 (.A1(n_2532_o_0),
    .A2(n_2551_o_0),
    .B(n_2557_o_0),
    .Y(n_2558_o_0));
 AOI21xp33_ASAP7_75t_R n_2559 (.A1(n_2394_o_0),
    .A2(n_2391_o_0),
    .B(ld),
    .Y(n_2559_o_0));
 AND2x2_ASAP7_75t_R n_2560 (.A(n_2415_o_0),
    .B(n_2543_o_0),
    .Y(n_2560_o_0));
 NAND2xp33_ASAP7_75t_R n_2561 (.A(net75),
    .B(n_2461_o_0),
    .Y(n_2561_o_0));
 NAND2xp33_ASAP7_75t_R n_2562 (.A(net75),
    .B(n_2506_o_0),
    .Y(n_2562_o_0));
 OAI21xp33_ASAP7_75t_R n_2563 (.A1(n_2498_o_0),
    .A2(net100),
    .B(net101),
    .Y(n_2563_o_0));
 AOI31xp67_ASAP7_75t_R n_2564 (.A1(n_2525_o_0),
    .A2(n_2523_o_0),
    .A3(n_827_o_0),
    .B(n_2526_o_0),
    .Y(n_2564_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2565 (.A1(n_2562_o_0),
    .A2(n_2563_o_0),
    .B(net52),
    .C(n_2564_o_0),
    .Y(n_2565_o_0));
 OAI21xp33_ASAP7_75t_R n_2566 (.A1(n_2498_o_0),
    .A2(net75),
    .B(n_2415_o_0),
    .Y(n_2566_o_0));
 NOR2xp33_ASAP7_75t_R n_2567 (.A(n_2498_o_0),
    .B(n_2484_o_0),
    .Y(n_2567_o_0));
 NAND2xp33_ASAP7_75t_R n_2568 (.A(n_2498_o_0),
    .B(n_2505_o_0),
    .Y(n_2568_o_0));
 INVx1_ASAP7_75t_R n_2569 (.A(n_2568_o_0),
    .Y(n_2569_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2570 (.A1(n_2567_o_0),
    .A2(n_2569_o_0),
    .B(n_2507_o_0),
    .C(n_2564_o_0),
    .Y(n_2570_o_0));
 OAI21xp33_ASAP7_75t_R n_2571 (.A1(n_2566_o_0),
    .A2(n_2540_o_0),
    .B(n_2570_o_0),
    .Y(n_2571_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2572 (.A1(n_2560_o_0),
    .A2(n_2561_o_0),
    .B(n_2565_o_0),
    .C(n_2571_o_0),
    .Y(n_2572_o_0));
 OAI221xp5_ASAP7_75t_R n_2573 (.A1(n_2437_o_0),
    .A2(n_2459_o_0),
    .B1(ld),
    .B2(n_2546_o_0),
    .C(n_2542_o_0),
    .Y(n_2573_o_0));
 NOR2xp33_ASAP7_75t_R n_2574 (.A(n_2437_o_0),
    .B(n_2459_o_0),
    .Y(n_2574_o_0));
 NAND2xp33_ASAP7_75t_R n_2575 (.A(n_2484_o_0),
    .B(n_2574_o_0),
    .Y(n_2575_o_0));
 NOR2xp33_ASAP7_75t_R n_2576 (.A(n_2498_o_0),
    .B(n_2459_o_0),
    .Y(n_2576_o_0));
 NOR3xp33_ASAP7_75t_R n_2577 (.A(n_2576_o_0),
    .B(n_2507_o_0),
    .C(net101),
    .Y(n_2577_o_0));
 AOI31xp33_ASAP7_75t_R n_2578 (.A1(n_2543_o_0),
    .A2(n_2575_o_0),
    .A3(n_2507_o_0),
    .B(n_2577_o_0),
    .Y(n_2578_o_0));
 OAI21xp33_ASAP7_75t_R n_2579 (.A1(n_2507_o_0),
    .A2(n_2573_o_0),
    .B(n_2578_o_0),
    .Y(n_2579_o_0));
 INVx1_ASAP7_75t_R n_2580 (.A(n_2546_o_0),
    .Y(n_2580_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2581 (.A1(n_2505_o_0),
    .A2(n_2498_o_0),
    .B(n_2538_o_0),
    .C(n_2542_o_0),
    .Y(n_2581_o_0));
 AOI211xp5_ASAP7_75t_R n_2582 (.A1(n_2580_o_0),
    .A2(n_827_o_0),
    .B(n_2581_o_0),
    .C(n_2507_o_0),
    .Y(n_2582_o_0));
 NOR2xp33_ASAP7_75t_R n_2583 (.A(net100),
    .B(n_2485_o_0),
    .Y(n_2583_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2584 (.A1(n_2539_o_0),
    .A2(n_827_o_0),
    .B(n_2504_o_0),
    .C(n_2437_o_0),
    .Y(n_2584_o_0));
 OAI21xp33_ASAP7_75t_R n_2585 (.A1(n_2459_o_0),
    .A2(n_2437_o_0),
    .B(n_2584_o_0),
    .Y(n_2585_o_0));
 AOI21xp33_ASAP7_75t_R n_2586 (.A1(net75),
    .A2(n_2585_o_0),
    .B(n_2415_o_0),
    .Y(n_2586_o_0));
 NOR4xp25_ASAP7_75t_R n_2587 (.A(n_2582_o_0),
    .B(n_2564_o_0),
    .C(n_2583_o_0),
    .D(n_2586_o_0),
    .Y(n_2587_o_0));
 AOI21xp33_ASAP7_75t_R n_2588 (.A1(n_2564_o_0),
    .A2(n_2579_o_0),
    .B(n_2587_o_0),
    .Y(n_2588_o_0));
 OAI321xp33_ASAP7_75t_R n_2589 (.A1(n_2559_o_0),
    .A2(n_2531_o_0),
    .A3(n_2572_o_0),
    .B1(n_2588_o_0),
    .B2(n_2532_o_0),
    .C(n_2385_o_0),
    .Y(n_2589_o_0));
 OAI31xp33_ASAP7_75t_R n_2590 (.A1(n_2385_o_0),
    .A2(n_2528_o_0),
    .A3(n_2558_o_0),
    .B(n_2589_o_0),
    .Y(n_2590_o_0));
 NAND2xp33_ASAP7_75t_R n_2591 (.A(n_2498_o_0),
    .B(n_2505_o_0),
    .Y(n_2591_o_0));
 AOI21xp33_ASAP7_75t_R n_2592 (.A1(n_2584_o_0),
    .A2(n_2591_o_0),
    .B(n_2492_o_0),
    .Y(n_2592_o_0));
 NOR2xp33_ASAP7_75t_R n_2593 (.A(net100),
    .B(net21),
    .Y(n_2593_o_0));
 AOI21xp33_ASAP7_75t_R n_2594 (.A1(n_2437_o_0),
    .A2(n_2492_o_0),
    .B(n_2415_o_0),
    .Y(n_2594_o_0));
 OAI21xp33_ASAP7_75t_R n_2595 (.A1(n_2576_o_0),
    .A2(net101),
    .B(n_2594_o_0),
    .Y(n_2595_o_0));
 OAI31xp33_ASAP7_75t_R n_2596 (.A1(n_2507_o_0),
    .A2(n_2592_o_0),
    .A3(n_2593_o_0),
    .B(n_2595_o_0),
    .Y(n_2596_o_0));
 INVx1_ASAP7_75t_R n_2597 (.A(n_2596_o_0),
    .Y(n_2597_o_0));
 OAI21xp33_ASAP7_75t_R n_2598 (.A1(n_2459_o_0),
    .A2(n_2437_o_0),
    .B(n_2484_o_0),
    .Y(n_2598_o_0));
 INVx1_ASAP7_75t_R n_2599 (.A(n_2598_o_0),
    .Y(n_2599_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2600 (.A1(n_2574_o_0),
    .A2(n_2492_o_0),
    .B(n_2599_o_0),
    .C(n_2415_o_0),
    .Y(n_2600_o_0));
 NAND3xp33_ASAP7_75t_R n_2601 (.A(n_2600_o_0),
    .B(n_2512_o_0),
    .C(n_2527_o_0),
    .Y(n_2601_o_0));
 OAI21xp33_ASAP7_75t_R n_2602 (.A1(n_2527_o_0),
    .A2(n_2597_o_0),
    .B(n_2601_o_0),
    .Y(n_2602_o_0));
 INVx1_ASAP7_75t_R n_2603 (.A(n_2559_o_0),
    .Y(n_2603_o_0));
 INVx1_ASAP7_75t_R n_2604 (.A(n_2531_o_0),
    .Y(n_2604_o_0));
 INVx1_ASAP7_75t_R n_2605 (.A(n_2543_o_0),
    .Y(n_2605_o_0));
 NAND3xp33_ASAP7_75t_R n_2606 (.A(n_2576_o_0),
    .B(n_2492_o_0),
    .C(n_2415_o_0),
    .Y(n_2606_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2607 (.A1(net52),
    .A2(n_2605_o_0),
    .B(n_2606_o_0),
    .C(n_2564_o_0),
    .Y(n_2607_o_0));
 NOR2xp33_ASAP7_75t_R n_2608 (.A(n_2415_o_0),
    .B(n_2484_o_0),
    .Y(n_2608_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2609 (.A1(n_2608_o_0),
    .A2(n_2460_o_0),
    .B(n_2499_o_0),
    .C(n_2564_o_0),
    .Y(n_2609_o_0));
 OAI21xp33_ASAP7_75t_R n_2610 (.A1(n_2510_o_0),
    .A2(n_2485_o_0),
    .B(n_2609_o_0),
    .Y(n_2610_o_0));
 AOI211xp5_ASAP7_75t_R n_2611 (.A1(n_2603_o_0),
    .A2(n_2604_o_0),
    .B(n_2607_o_0),
    .C(n_2610_o_0),
    .Y(n_2611_o_0));
 AOI21xp33_ASAP7_75t_R n_2612 (.A1(n_2602_o_0),
    .A2(n_2532_o_0),
    .B(n_2611_o_0),
    .Y(n_2612_o_0));
 OAI21xp33_ASAP7_75t_R n_2613 (.A1(n_2498_o_0),
    .A2(n_2492_o_0),
    .B(n_2415_o_0),
    .Y(n_2613_o_0));
 INVx1_ASAP7_75t_R n_2614 (.A(n_2613_o_0),
    .Y(n_2614_o_0));
 NOR3xp33_ASAP7_75t_R n_2615 (.A(n_2437_o_0),
    .B(n_2505_o_0),
    .C(n_2541_o_0),
    .Y(n_2615_o_0));
 OAI21xp33_ASAP7_75t_R n_2616 (.A1(n_2546_o_0),
    .A2(ld),
    .B(n_2615_o_0),
    .Y(n_2616_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2617 (.A1(n_2498_o_0),
    .A2(n_2492_o_0),
    .B(n_2573_o_0),
    .C(n_2415_o_0),
    .Y(n_2617_o_0));
 AO21x1_ASAP7_75t_R n_2618 (.A1(n_2614_o_0),
    .A2(n_2616_o_0),
    .B(n_2617_o_0),
    .Y(n_2618_o_0));
 NOR2xp33_ASAP7_75t_R n_2619 (.A(n_2505_o_0),
    .B(n_2484_o_0),
    .Y(n_2619_o_0));
 NAND2xp33_ASAP7_75t_R n_2620 (.A(n_2507_o_0),
    .B(n_2619_o_0),
    .Y(n_2620_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2621 (.A1(n_2585_o_0),
    .A2(n_2485_o_0),
    .B(n_2620_o_0),
    .C(n_2564_o_0),
    .Y(n_2621_o_0));
 AOI211xp5_ASAP7_75t_R n_2622 (.A1(n_2618_o_0),
    .A2(n_2564_o_0),
    .B(n_2532_o_0),
    .C(n_2621_o_0),
    .Y(n_2622_o_0));
 AOI21xp33_ASAP7_75t_R n_2623 (.A1(net21),
    .A2(n_2576_o_0),
    .B(n_2507_o_0),
    .Y(n_2623_o_0));
 OAI31xp33_ASAP7_75t_R n_2624 (.A1(net52),
    .A2(n_2506_o_0),
    .A3(net21),
    .B(n_2527_o_0),
    .Y(n_2624_o_0));
 OAI221xp5_ASAP7_75t_R n_2625 (.A1(n_2498_o_0),
    .A2(net100),
    .B1(ld),
    .B2(n_2580_o_0),
    .C(n_2482_o_0),
    .Y(n_2625_o_0));
 AOI311xp33_ASAP7_75t_R n_2626 (.A1(n_2507_o_0),
    .A2(n_2616_o_0),
    .A3(n_2625_o_0),
    .B(n_2527_o_0),
    .C(n_2508_o_0),
    .Y(n_2626_o_0));
 INVx1_ASAP7_75t_R n_2627 (.A(n_2626_o_0),
    .Y(n_2627_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2628 (.A1(n_2616_o_0),
    .A2(n_2623_o_0),
    .B(n_2624_o_0),
    .C(n_2627_o_0),
    .D(n_2396_o_0),
    .Y(n_2628_o_0));
 OAI31xp33_ASAP7_75t_R n_2629 (.A1(n_2622_o_0),
    .A2(n_2628_o_0),
    .A3(n_2384_o_0),
    .B(n_2372_o_0),
    .Y(n_2629_o_0));
 AOI21xp33_ASAP7_75t_R n_2630 (.A1(n_2384_o_0),
    .A2(n_2612_o_0),
    .B(n_2629_o_0),
    .Y(n_2630_o_0));
 AOI21xp33_ASAP7_75t_R n_2631 (.A1(n_2373_o_0),
    .A2(n_2590_o_0),
    .B(n_2630_o_0),
    .Y(n_2631_o_0));
 NAND2xp33_ASAP7_75t_R n_2632 (.A(n_2492_o_0),
    .B(n_2460_o_0),
    .Y(n_2632_o_0));
 AOI21xp33_ASAP7_75t_R n_2633 (.A1(n_2498_o_0),
    .A2(net100),
    .B(n_2541_o_0),
    .Y(n_2633_o_0));
 OAI21xp33_ASAP7_75t_R n_2634 (.A1(n_2546_o_0),
    .A2(ld),
    .B(n_2633_o_0),
    .Y(n_2634_o_0));
 INVx1_ASAP7_75t_R n_2635 (.A(n_2634_o_0),
    .Y(n_2635_o_0));
 AOI22xp33_ASAP7_75t_R n_2636 (.A1(n_2586_o_0),
    .A2(n_2632_o_0),
    .B1(net52),
    .B2(n_2635_o_0),
    .Y(n_2636_o_0));
 NOR2xp33_ASAP7_75t_R n_2637 (.A(n_2505_o_0),
    .B(net101),
    .Y(n_2637_o_0));
 AOI21xp33_ASAP7_75t_R n_2638 (.A1(n_2507_o_0),
    .A2(n_2637_o_0),
    .B(n_2564_o_0),
    .Y(n_2638_o_0));
 OAI21xp33_ASAP7_75t_R n_2639 (.A1(n_2510_o_0),
    .A2(n_2485_o_0),
    .B(n_2396_o_0),
    .Y(n_2639_o_0));
 AOI21xp33_ASAP7_75t_R n_2640 (.A1(n_2554_o_0),
    .A2(n_2638_o_0),
    .B(n_2639_o_0),
    .Y(n_2640_o_0));
 OAI21xp33_ASAP7_75t_R n_2641 (.A1(n_2527_o_0),
    .A2(n_2636_o_0),
    .B(n_2640_o_0),
    .Y(n_2641_o_0));
 NAND2xp33_ASAP7_75t_R n_2642 (.A(net102),
    .B(net75),
    .Y(n_2642_o_0));
 INVx1_ASAP7_75t_R n_2643 (.A(n_2642_o_0),
    .Y(n_2643_o_0));
 NAND2xp33_ASAP7_75t_R n_2644 (.A(n_2492_o_0),
    .B(n_2510_o_0),
    .Y(n_2644_o_0));
 INVx1_ASAP7_75t_R n_2645 (.A(n_2644_o_0),
    .Y(n_2645_o_0));
 NAND3xp33_ASAP7_75t_R n_2646 (.A(n_2543_o_0),
    .B(n_2552_o_0),
    .C(n_2507_o_0),
    .Y(n_2646_o_0));
 OAI31xp33_ASAP7_75t_R n_2647 (.A1(n_2507_o_0),
    .A2(n_2643_o_0),
    .A3(n_2645_o_0),
    .B(n_2646_o_0),
    .Y(n_2647_o_0));
 NAND2xp33_ASAP7_75t_R n_2648 (.A(n_2459_o_0),
    .B(n_2492_o_0),
    .Y(n_2648_o_0));
 AOI211xp5_ASAP7_75t_R n_2649 (.A1(net100),
    .A2(n_2498_o_0),
    .B(net101),
    .C(n_2415_o_0),
    .Y(n_2649_o_0));
 AOI31xp33_ASAP7_75t_R n_2650 (.A1(net52),
    .A2(n_2568_o_0),
    .A3(n_2648_o_0),
    .B(n_2649_o_0),
    .Y(n_2650_o_0));
 OAI21xp33_ASAP7_75t_R n_2651 (.A1(n_2527_o_0),
    .A2(n_2650_o_0),
    .B(n_2532_o_0),
    .Y(n_2651_o_0));
 AO21x1_ASAP7_75t_R n_2652 (.A1(n_2647_o_0),
    .A2(n_2527_o_0),
    .B(n_2651_o_0),
    .Y(n_2652_o_0));
 AOI211xp5_ASAP7_75t_R n_2653 (.A1(net100),
    .A2(n_2437_o_0),
    .B(n_2507_o_0),
    .C(net75),
    .Y(n_2653_o_0));
 AOI21xp33_ASAP7_75t_R n_2654 (.A1(n_2505_o_0),
    .A2(n_2492_o_0),
    .B(n_2415_o_0),
    .Y(n_2654_o_0));
 OAI211xp5_ASAP7_75t_R n_2655 (.A1(n_2653_o_0),
    .A2(n_2654_o_0),
    .B(n_2545_o_0),
    .C(n_2527_o_0),
    .Y(n_2655_o_0));
 AOI211xp5_ASAP7_75t_R n_2656 (.A1(key[26]),
    .A2(ld),
    .B(n_2505_o_0),
    .C(n_2498_o_0),
    .Y(n_2656_o_0));
 OAI21xp33_ASAP7_75t_R n_2657 (.A1(ld),
    .A2(n_2580_o_0),
    .B(n_2656_o_0),
    .Y(n_2657_o_0));
 OAI211xp5_ASAP7_75t_R n_2658 (.A1(n_2585_o_0),
    .A2(net75),
    .B(n_2657_o_0),
    .C(n_2507_o_0),
    .Y(n_2658_o_0));
 OAI31xp33_ASAP7_75t_R n_2659 (.A1(n_2507_o_0),
    .A2(net21),
    .A3(n_2510_o_0),
    .B(n_2658_o_0),
    .Y(n_2659_o_0));
 AOI21xp33_ASAP7_75t_R n_2660 (.A1(n_2564_o_0),
    .A2(n_2659_o_0),
    .B(n_2396_o_0),
    .Y(n_2660_o_0));
 INVx1_ASAP7_75t_R n_2661 (.A(n_2573_o_0),
    .Y(n_2661_o_0));
 OAI211xp5_ASAP7_75t_R n_2662 (.A1(n_2546_o_0),
    .A2(ld),
    .B(n_2585_o_0),
    .C(n_2542_o_0),
    .Y(n_2662_o_0));
 AOI21xp33_ASAP7_75t_R n_2663 (.A1(net21),
    .A2(n_2511_o_0),
    .B(n_2415_o_0),
    .Y(n_2663_o_0));
 AOI21xp33_ASAP7_75t_R n_2664 (.A1(n_2662_o_0),
    .A2(n_2663_o_0),
    .B(n_2564_o_0),
    .Y(n_2664_o_0));
 INVx1_ASAP7_75t_R n_2665 (.A(n_2592_o_0),
    .Y(n_2665_o_0));
 OAI21xp33_ASAP7_75t_R n_2666 (.A1(n_2498_o_0),
    .A2(n_2484_o_0),
    .B(n_2415_o_0),
    .Y(n_2666_o_0));
 INVx1_ASAP7_75t_R n_2667 (.A(n_2666_o_0),
    .Y(n_2667_o_0));
 OAI21xp33_ASAP7_75t_R n_2668 (.A1(n_2437_o_0),
    .A2(n_2484_o_0),
    .B(n_2507_o_0),
    .Y(n_2668_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2669 (.A1(net100),
    .A2(net102),
    .B(n_2668_o_0),
    .C(n_2564_o_0),
    .Y(n_2669_o_0));
 AOI21xp33_ASAP7_75t_R n_2670 (.A1(n_2665_o_0),
    .A2(n_2667_o_0),
    .B(n_2669_o_0),
    .Y(n_2670_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2671 (.A1(n_2661_o_0),
    .A2(n_2613_o_0),
    .B(n_2664_o_0),
    .C(n_2670_o_0),
    .Y(n_2671_o_0));
 AOI221xp5_ASAP7_75t_R n_2672 (.A1(n_2655_o_0),
    .A2(n_2660_o_0),
    .B1(n_2396_o_0),
    .B2(n_2671_o_0),
    .C(n_2385_o_0),
    .Y(n_2672_o_0));
 AOI31xp33_ASAP7_75t_R n_2673 (.A1(n_2385_o_0),
    .A2(n_2641_o_0),
    .A3(n_2652_o_0),
    .B(n_2672_o_0),
    .Y(n_2673_o_0));
 NAND2xp33_ASAP7_75t_R n_2674 (.A(n_2459_o_0),
    .B(n_2484_o_0),
    .Y(n_2674_o_0));
 INVx1_ASAP7_75t_R n_2675 (.A(n_2674_o_0),
    .Y(n_2675_o_0));
 NOR2xp33_ASAP7_75t_R n_2676 (.A(n_2666_o_0),
    .B(n_2675_o_0),
    .Y(n_2676_o_0));
 NOR2xp33_ASAP7_75t_R n_2677 (.A(n_2459_o_0),
    .B(n_2492_o_0),
    .Y(n_2677_o_0));
 NOR2xp33_ASAP7_75t_R n_2678 (.A(n_2677_o_0),
    .B(n_2512_o_0),
    .Y(n_2678_o_0));
 OAI21xp33_ASAP7_75t_R n_2679 (.A1(n_2676_o_0),
    .A2(n_2678_o_0),
    .B(n_2396_o_0),
    .Y(n_2679_o_0));
 AOI21xp33_ASAP7_75t_R n_2680 (.A1(n_2492_o_0),
    .A2(n_2498_o_0),
    .B(n_2507_o_0),
    .Y(n_2680_o_0));
 AOI21xp33_ASAP7_75t_R n_2681 (.A1(n_2680_o_0),
    .A2(n_2575_o_0),
    .B(n_2649_o_0),
    .Y(n_2681_o_0));
 OAI21xp33_ASAP7_75t_R n_2682 (.A1(net52),
    .A2(n_2632_o_0),
    .B(n_2681_o_0),
    .Y(n_2682_o_0));
 AOI21xp33_ASAP7_75t_R n_2683 (.A1(n_2532_o_0),
    .A2(n_2682_o_0),
    .B(n_2564_o_0),
    .Y(n_2683_o_0));
 NAND2xp33_ASAP7_75t_R n_2684 (.A(n_2505_o_0),
    .B(net75),
    .Y(n_2684_o_0));
 AOI31xp33_ASAP7_75t_R n_2685 (.A1(n_2459_o_0),
    .A2(n_2437_o_0),
    .A3(n_2492_o_0),
    .B(n_2507_o_0),
    .Y(n_2685_o_0));
 NAND3xp33_ASAP7_75t_R n_2686 (.A(net75),
    .B(n_2437_o_0),
    .C(n_2505_o_0),
    .Y(n_2686_o_0));
 AOI32xp33_ASAP7_75t_R n_2687 (.A1(n_2684_o_0),
    .A2(n_2396_o_0),
    .A3(n_2507_o_0),
    .B1(n_2685_o_0),
    .B2(n_2686_o_0),
    .Y(n_2687_o_0));
 AO21x1_ASAP7_75t_R n_2688 (.A1(n_2687_o_0),
    .A2(n_2564_o_0),
    .B(n_2384_o_0),
    .Y(n_2688_o_0));
 AOI21xp33_ASAP7_75t_R n_2689 (.A1(n_2679_o_0),
    .A2(n_2683_o_0),
    .B(n_2688_o_0),
    .Y(n_2689_o_0));
 NAND2xp33_ASAP7_75t_R n_2690 (.A(n_2505_o_0),
    .B(n_2484_o_0),
    .Y(n_2690_o_0));
 INVx1_ASAP7_75t_R n_2691 (.A(n_2690_o_0),
    .Y(n_2691_o_0));
 NAND2xp33_ASAP7_75t_R n_2692 (.A(n_2575_o_0),
    .B(n_2667_o_0),
    .Y(n_2692_o_0));
 OAI31xp33_ASAP7_75t_R n_2693 (.A1(n_2645_o_0),
    .A2(n_2691_o_0),
    .A3(net52),
    .B(n_2692_o_0),
    .Y(n_2693_o_0));
 AOI21xp33_ASAP7_75t_R n_2694 (.A1(n_2507_o_0),
    .A2(n_2543_o_0),
    .B(n_2653_o_0),
    .Y(n_2694_o_0));
 NAND2xp33_ASAP7_75t_R n_2695 (.A(net102),
    .B(net75),
    .Y(n_2695_o_0));
 AOI31xp33_ASAP7_75t_R n_2696 (.A1(n_2396_o_0),
    .A2(n_2694_o_0),
    .A3(n_2695_o_0),
    .B(n_2527_o_0),
    .Y(n_2696_o_0));
 OAI21xp33_ASAP7_75t_R n_2697 (.A1(n_2396_o_0),
    .A2(n_2693_o_0),
    .B(n_2696_o_0),
    .Y(n_2697_o_0));
 AOI21xp33_ASAP7_75t_R n_2698 (.A1(n_2492_o_0),
    .A2(n_2460_o_0),
    .B(n_2507_o_0),
    .Y(n_2698_o_0));
 NOR2xp33_ASAP7_75t_R n_2699 (.A(net21),
    .B(n_2585_o_0),
    .Y(n_2699_o_0));
 NAND2xp33_ASAP7_75t_R n_2700 (.A(n_2507_o_0),
    .B(n_2657_o_0),
    .Y(n_2700_o_0));
 OAI21xp33_ASAP7_75t_R n_2701 (.A1(n_2699_o_0),
    .A2(n_2700_o_0),
    .B(n_2396_o_0),
    .Y(n_2701_o_0));
 NAND2xp33_ASAP7_75t_R n_2702 (.A(n_2484_o_0),
    .B(n_2507_o_0),
    .Y(n_2702_o_0));
 OA222x2_ASAP7_75t_R n_2703 (.A1(n_2585_o_0),
    .A2(n_2702_o_0),
    .B1(n_2573_o_0),
    .B2(n_2415_o_0),
    .C1(n_2485_o_0),
    .C2(n_2498_o_0),
    .Y(n_2703_o_0));
 INVx1_ASAP7_75t_R n_2704 (.A(n_2508_o_0),
    .Y(n_2704_o_0));
 AOI31xp33_ASAP7_75t_R n_2705 (.A1(n_2532_o_0),
    .A2(n_2703_o_0),
    .A3(n_2704_o_0),
    .B(n_2564_o_0),
    .Y(n_2705_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2706 (.A1(n_2598_o_0),
    .A2(n_2698_o_0),
    .B(n_2701_o_0),
    .C(n_2705_o_0),
    .Y(n_2706_o_0));
 AOI21xp33_ASAP7_75t_R n_2707 (.A1(n_2697_o_0),
    .A2(n_2706_o_0),
    .B(n_2385_o_0),
    .Y(n_2707_o_0));
 OAI21xp33_ASAP7_75t_R n_2708 (.A1(n_2689_o_0),
    .A2(n_2707_o_0),
    .B(n_2373_o_0),
    .Y(n_2708_o_0));
 OAI21xp33_ASAP7_75t_R n_2709 (.A1(n_2373_o_0),
    .A2(n_2673_o_0),
    .B(n_2708_o_0),
    .Y(n_2709_o_0));
 NAND2xp33_ASAP7_75t_R n_2710 (.A(n_2484_o_0),
    .B(n_2510_o_0),
    .Y(n_2710_o_0));
 AOI21xp33_ASAP7_75t_R n_2711 (.A1(n_2710_o_0),
    .A2(n_2544_o_0),
    .B(n_2527_o_0),
    .Y(n_2711_o_0));
 AO21x1_ASAP7_75t_R n_2712 (.A1(n_2685_o_0),
    .A2(n_2686_o_0),
    .B(n_2564_o_0),
    .Y(n_2712_o_0));
 AOI21xp33_ASAP7_75t_R n_2713 (.A1(n_2594_o_0),
    .A2(n_2657_o_0),
    .B(n_2712_o_0),
    .Y(n_2713_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2714 (.A1(n_2507_o_0),
    .A2(n_2573_o_0),
    .B(n_2711_o_0),
    .C(n_2713_o_0),
    .Y(n_2714_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2715 (.A1(n_827_o_0),
    .A2(n_2546_o_0),
    .B(n_2547_o_0),
    .C(n_2415_o_0),
    .Y(n_2715_o_0));
 OAI21xp33_ASAP7_75t_R n_2716 (.A1(n_2619_o_0),
    .A2(n_2415_o_0),
    .B(n_2715_o_0),
    .Y(n_2716_o_0));
 INVx1_ASAP7_75t_R n_2717 (.A(n_2716_o_0),
    .Y(n_2717_o_0));
 INVx1_ASAP7_75t_R n_2718 (.A(n_2648_o_0),
    .Y(n_2718_o_0));
 OAI31xp33_ASAP7_75t_R n_2719 (.A1(net52),
    .A2(n_2718_o_0),
    .A3(n_2555_o_0),
    .B(n_2527_o_0),
    .Y(n_2719_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2720 (.A1(net52),
    .A2(n_2637_o_0),
    .B(n_2719_o_0),
    .C(n_2396_o_0),
    .Y(n_2720_o_0));
 AOI21xp33_ASAP7_75t_R n_2721 (.A1(n_2717_o_0),
    .A2(n_2564_o_0),
    .B(n_2720_o_0),
    .Y(n_2721_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2722 (.A1(n_2714_o_0),
    .A2(n_2532_o_0),
    .B(n_2721_o_0),
    .C(n_2372_o_0),
    .Y(n_2722_o_0));
 NAND2xp33_ASAP7_75t_R n_2723 (.A(n_2594_o_0),
    .B(n_2575_o_0),
    .Y(n_2723_o_0));
 OAI31xp33_ASAP7_75t_R n_2724 (.A1(n_2507_o_0),
    .A2(n_2699_o_0),
    .A3(n_2691_o_0),
    .B(n_2723_o_0),
    .Y(n_2724_o_0));
 NAND2xp33_ASAP7_75t_R n_2725 (.A(n_2564_o_0),
    .B(n_2715_o_0),
    .Y(n_2725_o_0));
 AOI31xp33_ASAP7_75t_R n_2726 (.A1(n_2657_o_0),
    .A2(n_2507_o_0),
    .A3(n_2632_o_0),
    .B(n_2725_o_0),
    .Y(n_2726_o_0));
 AOI21xp33_ASAP7_75t_R n_2727 (.A1(n_2527_o_0),
    .A2(n_2724_o_0),
    .B(n_2726_o_0),
    .Y(n_2727_o_0));
 NOR3xp33_ASAP7_75t_R n_2728 (.A(n_2718_o_0),
    .B(n_2555_o_0),
    .C(n_2415_o_0),
    .Y(n_2728_o_0));
 AOI31xp33_ASAP7_75t_R n_2729 (.A1(net52),
    .A2(n_2545_o_0),
    .A3(n_2644_o_0),
    .B(n_2728_o_0),
    .Y(n_2729_o_0));
 NOR3xp33_ASAP7_75t_R n_2730 (.A(n_2452_o_0),
    .B(n_2457_o_0),
    .C(ld),
    .Y(n_2730_o_0));
 NOR2xp33_ASAP7_75t_R n_2731 (.A(n_2534_o_0),
    .B(n_827_o_0),
    .Y(n_2731_o_0));
 OAI311xp33_ASAP7_75t_R n_2732 (.A1(n_2730_o_0),
    .A2(n_2731_o_0),
    .A3(n_2437_o_0),
    .B1(n_2484_o_0),
    .C1(n_2584_o_0),
    .Y(n_2732_o_0));
 INVx1_ASAP7_75t_R n_2733 (.A(n_2732_o_0),
    .Y(n_2733_o_0));
 AOI21xp33_ASAP7_75t_R n_2734 (.A1(n_2459_o_0),
    .A2(n_2492_o_0),
    .B(n_2507_o_0),
    .Y(n_2734_o_0));
 INVx1_ASAP7_75t_R n_2735 (.A(n_2734_o_0),
    .Y(n_2735_o_0));
 AOI21xp33_ASAP7_75t_R n_2736 (.A1(n_2634_o_0),
    .A2(n_2663_o_0),
    .B(n_2527_o_0),
    .Y(n_2736_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2737 (.A1(n_2733_o_0),
    .A2(n_2735_o_0),
    .B(n_2736_o_0),
    .C(n_2532_o_0),
    .Y(n_2737_o_0));
 OAI21xp33_ASAP7_75t_R n_2738 (.A1(n_2564_o_0),
    .A2(n_2729_o_0),
    .B(n_2737_o_0),
    .Y(n_2738_o_0));
 OAI211xp5_ASAP7_75t_R n_2739 (.A1(n_2396_o_0),
    .A2(n_2727_o_0),
    .B(n_2738_o_0),
    .C(n_2373_o_0),
    .Y(n_2739_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2740 (.A1(net102),
    .A2(net21),
    .B(n_2505_o_0),
    .C(net52),
    .Y(n_2740_o_0));
 OAI21xp33_ASAP7_75t_R n_2741 (.A1(n_2492_o_0),
    .A2(n_2460_o_0),
    .B(n_2415_o_0),
    .Y(n_2741_o_0));
 OAI21xp33_ASAP7_75t_R n_2742 (.A1(n_2567_o_0),
    .A2(n_2741_o_0),
    .B(n_2527_o_0),
    .Y(n_2742_o_0));
 NOR2xp33_ASAP7_75t_R n_2743 (.A(net101),
    .B(n_2585_o_0),
    .Y(n_2743_o_0));
 INVx1_ASAP7_75t_R n_2744 (.A(n_2743_o_0),
    .Y(n_2744_o_0));
 OAI221xp5_ASAP7_75t_R n_2745 (.A1(n_2498_o_0),
    .A2(n_2459_o_0),
    .B1(ld),
    .B2(n_2580_o_0),
    .C(n_2482_o_0),
    .Y(n_2745_o_0));
 INVx1_ASAP7_75t_R n_2746 (.A(n_2745_o_0),
    .Y(n_2746_o_0));
 AOI211xp5_ASAP7_75t_R n_2747 (.A1(net101),
    .A2(n_2498_o_0),
    .B(n_2746_o_0),
    .C(n_2507_o_0),
    .Y(n_2747_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2748 (.A1(n_2544_o_0),
    .A2(n_2744_o_0),
    .B(n_2747_o_0),
    .C(n_2564_o_0),
    .Y(n_2748_o_0));
 OAI211xp5_ASAP7_75t_R n_2749 (.A1(n_2740_o_0),
    .A2(n_2742_o_0),
    .B(n_2748_o_0),
    .C(n_2532_o_0),
    .Y(n_2749_o_0));
 INVx1_ASAP7_75t_R n_2750 (.A(n_2654_o_0),
    .Y(n_2750_o_0));
 AOI21xp33_ASAP7_75t_R n_2751 (.A1(n_2510_o_0),
    .A2(net21),
    .B(n_2750_o_0),
    .Y(n_2751_o_0));
 OAI21xp33_ASAP7_75t_R n_2752 (.A1(n_2510_o_0),
    .A2(n_2485_o_0),
    .B(n_2606_o_0),
    .Y(n_2752_o_0));
 OAI21xp33_ASAP7_75t_R n_2753 (.A1(net101),
    .A2(n_2510_o_0),
    .B(n_2507_o_0),
    .Y(n_2753_o_0));
 OAI21xp33_ASAP7_75t_R n_2754 (.A1(n_2567_o_0),
    .A2(n_2753_o_0),
    .B(n_2741_o_0),
    .Y(n_2754_o_0));
 NAND3xp33_ASAP7_75t_R n_2755 (.A(n_2754_o_0),
    .B(n_2606_o_0),
    .C(n_2527_o_0),
    .Y(n_2755_o_0));
 OAI31xp33_ASAP7_75t_R n_2756 (.A1(n_2527_o_0),
    .A2(n_2751_o_0),
    .A3(n_2752_o_0),
    .B(n_2755_o_0),
    .Y(n_2756_o_0));
 AOI21xp33_ASAP7_75t_R n_2757 (.A1(n_2396_o_0),
    .A2(n_2756_o_0),
    .B(n_2372_o_0),
    .Y(n_2757_o_0));
 AOI21xp33_ASAP7_75t_R n_2758 (.A1(n_2749_o_0),
    .A2(n_2757_o_0),
    .B(n_2385_o_0),
    .Y(n_2758_o_0));
 NOR2xp33_ASAP7_75t_R n_2759 (.A(n_2668_o_0),
    .B(n_2691_o_0),
    .Y(n_2759_o_0));
 AOI31xp33_ASAP7_75t_R n_2760 (.A1(net52),
    .A2(n_2744_o_0),
    .A3(n_2648_o_0),
    .B(n_2759_o_0),
    .Y(n_2760_o_0));
 AOI21xp33_ASAP7_75t_R n_2761 (.A1(n_2532_o_0),
    .A2(n_2760_o_0),
    .B(n_2564_o_0),
    .Y(n_2761_o_0));
 AOI22xp33_ASAP7_75t_R n_2762 (.A1(n_2586_o_0),
    .A2(n_2616_o_0),
    .B1(net52),
    .B2(n_2619_o_0),
    .Y(n_2762_o_0));
 AOI21xp33_ASAP7_75t_R n_2763 (.A1(n_2532_o_0),
    .A2(n_2762_o_0),
    .B(n_2527_o_0),
    .Y(n_2763_o_0));
 NAND3xp33_ASAP7_75t_R n_2764 (.A(n_2648_o_0),
    .B(n_2568_o_0),
    .C(n_2507_o_0),
    .Y(n_2764_o_0));
 INVx1_ASAP7_75t_R n_2765 (.A(n_2764_o_0),
    .Y(n_2765_o_0));
 AOI21xp33_ASAP7_75t_R n_2766 (.A1(net52),
    .A2(n_2684_o_0),
    .B(n_2765_o_0),
    .Y(n_2766_o_0));
 NAND3xp33_ASAP7_75t_R n_2767 (.A(n_2732_o_0),
    .B(n_2563_o_0),
    .C(n_2507_o_0),
    .Y(n_2767_o_0));
 AOI21xp33_ASAP7_75t_R n_2768 (.A1(n_2734_o_0),
    .A2(n_2562_o_0),
    .B(n_2564_o_0),
    .Y(n_2768_o_0));
 AOI21xp33_ASAP7_75t_R n_2769 (.A1(n_2767_o_0),
    .A2(n_2768_o_0),
    .B(n_2532_o_0),
    .Y(n_2769_o_0));
 OAI21xp33_ASAP7_75t_R n_2770 (.A1(n_2527_o_0),
    .A2(n_2766_o_0),
    .B(n_2769_o_0),
    .Y(n_2770_o_0));
 OAI211xp5_ASAP7_75t_R n_2771 (.A1(n_2761_o_0),
    .A2(n_2763_o_0),
    .B(n_2770_o_0),
    .C(n_2372_o_0),
    .Y(n_2771_o_0));
 AOI32xp33_ASAP7_75t_R n_2772 (.A1(n_2722_o_0),
    .A2(n_2739_o_0),
    .A3(n_2385_o_0),
    .B1(n_2758_o_0),
    .B2(n_2771_o_0),
    .Y(n_2772_o_0));
 INVx1_ASAP7_75t_R n_2773 (.A(n_2576_o_0),
    .Y(n_2773_o_0));
 NAND2xp33_ASAP7_75t_R n_2774 (.A(net75),
    .B(n_2773_o_0),
    .Y(n_2774_o_0));
 INVx1_ASAP7_75t_R n_2775 (.A(n_2570_o_0),
    .Y(n_2775_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2776 (.A1(n_2591_o_0),
    .A2(n_2584_o_0),
    .B(net101),
    .C(n_2685_o_0),
    .Y(n_2776_o_0));
 OAI31xp33_ASAP7_75t_R n_2777 (.A1(net21),
    .A2(n_2576_o_0),
    .A3(net52),
    .B(n_2776_o_0),
    .Y(n_2777_o_0));
 OAI21xp33_ASAP7_75t_R n_2778 (.A1(n_2649_o_0),
    .A2(n_2777_o_0),
    .B(n_2564_o_0),
    .Y(n_2778_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2779 (.A1(n_2774_o_0),
    .A2(n_2560_o_0),
    .B(n_2775_o_0),
    .C(n_2778_o_0),
    .D(n_2396_o_0),
    .Y(n_2779_o_0));
 AOI21xp33_ASAP7_75t_R n_2780 (.A1(n_2591_o_0),
    .A2(n_2695_o_0),
    .B(n_2507_o_0),
    .Y(n_2780_o_0));
 OAI21xp33_ASAP7_75t_R n_2781 (.A1(net52),
    .A2(n_2555_o_0),
    .B(n_2564_o_0),
    .Y(n_2781_o_0));
 INVx1_ASAP7_75t_R n_2782 (.A(n_2545_o_0),
    .Y(n_2782_o_0));
 AOI31xp33_ASAP7_75t_R n_2783 (.A1(n_2492_o_0),
    .A2(n_2591_o_0),
    .A3(n_2584_o_0),
    .B(n_2507_o_0),
    .Y(n_2783_o_0));
 AOI21xp33_ASAP7_75t_R n_2784 (.A1(n_2745_o_0),
    .A2(n_2783_o_0),
    .B(n_2564_o_0),
    .Y(n_2784_o_0));
 OAI21xp33_ASAP7_75t_R n_2785 (.A1(n_2782_o_0),
    .A2(n_2750_o_0),
    .B(n_2784_o_0),
    .Y(n_2785_o_0));
 OAI21xp33_ASAP7_75t_R n_2786 (.A1(n_2780_o_0),
    .A2(n_2781_o_0),
    .B(n_2785_o_0),
    .Y(n_2786_o_0));
 OAI21xp33_ASAP7_75t_R n_2787 (.A1(n_2532_o_0),
    .A2(n_2786_o_0),
    .B(n_2384_o_0),
    .Y(n_2787_o_0));
 AOI22xp33_ASAP7_75t_R n_2788 (.A1(n_2586_o_0),
    .A2(n_2573_o_0),
    .B1(n_2563_o_0),
    .B2(n_2614_o_0),
    .Y(n_2788_o_0));
 INVx1_ASAP7_75t_R n_2789 (.A(n_2553_o_0),
    .Y(n_2789_o_0));
 AOI21xp33_ASAP7_75t_R n_2790 (.A1(n_2690_o_0),
    .A2(n_2783_o_0),
    .B(n_2527_o_0),
    .Y(n_2790_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2791 (.A1(n_2510_o_0),
    .A2(net21),
    .B(n_2789_o_0),
    .C(n_2790_o_0),
    .Y(n_2791_o_0));
 OAI21xp33_ASAP7_75t_R n_2792 (.A1(n_2564_o_0),
    .A2(n_2788_o_0),
    .B(n_2791_o_0),
    .Y(n_2792_o_0));
 NOR2xp33_ASAP7_75t_R n_2793 (.A(n_2415_o_0),
    .B(n_2492_o_0),
    .Y(n_2793_o_0));
 AO21x1_ASAP7_75t_R n_2794 (.A1(n_2585_o_0),
    .A2(n_2793_o_0),
    .B(n_2564_o_0),
    .Y(n_2794_o_0));
 OAI21xp33_ASAP7_75t_R n_2795 (.A1(n_2794_o_0),
    .A2(n_2676_o_0),
    .B(n_2396_o_0),
    .Y(n_2795_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2796 (.A1(n_2690_o_0),
    .A2(n_2544_o_0),
    .B(n_2780_o_0),
    .C(n_2564_o_0),
    .D(n_2795_o_0),
    .Y(n_2796_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2797 (.A1(n_2532_o_0),
    .A2(n_2792_o_0),
    .B(n_2796_o_0),
    .C(n_2385_o_0),
    .Y(n_2797_o_0));
 OAI21xp33_ASAP7_75t_R n_2798 (.A1(n_2779_o_0),
    .A2(n_2787_o_0),
    .B(n_2797_o_0),
    .Y(n_2798_o_0));
 AOI22xp33_ASAP7_75t_R n_2799 (.A1(n_2585_o_0),
    .A2(n_2793_o_0),
    .B1(n_2686_o_0),
    .B2(n_2648_o_0),
    .Y(n_2799_o_0));
 NAND3xp33_ASAP7_75t_R n_2800 (.A(n_2585_o_0),
    .B(net21),
    .C(n_2507_o_0),
    .Y(n_2800_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2801 (.A1(n_2507_o_0),
    .A2(n_2799_o_0),
    .B(n_2800_o_0),
    .C(n_2532_o_0),
    .Y(n_2801_o_0));
 AOI31xp33_ASAP7_75t_R n_2802 (.A1(net101),
    .A2(n_2574_o_0),
    .A3(n_2507_o_0),
    .B(n_2801_o_0),
    .Y(n_2802_o_0));
 AOI21xp33_ASAP7_75t_R n_2803 (.A1(n_2532_o_0),
    .A2(n_2582_o_0),
    .B(n_2564_o_0),
    .Y(n_2803_o_0));
 NOR2xp33_ASAP7_75t_R n_2804 (.A(n_2415_o_0),
    .B(net75),
    .Y(n_2804_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2805 (.A1(n_2804_o_0),
    .A2(n_2576_o_0),
    .B(n_2747_o_0),
    .C(n_2532_o_0),
    .Y(n_2805_o_0));
 INVx1_ASAP7_75t_R n_2806 (.A(n_2594_o_0),
    .Y(n_2806_o_0));
 OAI211xp5_ASAP7_75t_R n_2807 (.A1(net102),
    .A2(net101),
    .B(n_2543_o_0),
    .C(n_2415_o_0),
    .Y(n_2807_o_0));
 OAI21xp33_ASAP7_75t_R n_2808 (.A1(n_2782_o_0),
    .A2(n_2806_o_0),
    .B(n_2807_o_0),
    .Y(n_2808_o_0));
 AOI21xp33_ASAP7_75t_R n_2809 (.A1(n_2396_o_0),
    .A2(n_2808_o_0),
    .B(n_2527_o_0),
    .Y(n_2809_o_0));
 AOI22xp33_ASAP7_75t_R n_2810 (.A1(n_2802_o_0),
    .A2(n_2803_o_0),
    .B1(n_2805_o_0),
    .B2(n_2809_o_0),
    .Y(n_2810_o_0));
 AOI22xp33_ASAP7_75t_R n_2811 (.A1(n_2685_o_0),
    .A2(n_2686_o_0),
    .B1(n_2594_o_0),
    .B2(n_2745_o_0),
    .Y(n_2811_o_0));
 OA21x2_ASAP7_75t_R n_2812 (.A1(n_2811_o_0),
    .A2(n_2527_o_0),
    .B(n_2396_o_0),
    .Y(n_2812_o_0));
 NOR2xp33_ASAP7_75t_R n_2813 (.A(net101),
    .B(n_2461_o_0),
    .Y(n_2813_o_0));
 AOI32xp33_ASAP7_75t_R n_2814 (.A1(n_2507_o_0),
    .A2(n_2498_o_0),
    .A3(net21),
    .B1(n_2608_o_0),
    .B2(n_2576_o_0),
    .Y(n_2814_o_0));
 OAI31xp33_ASAP7_75t_R n_2815 (.A1(n_2507_o_0),
    .A2(n_2605_o_0),
    .A3(n_2813_o_0),
    .B(n_2814_o_0),
    .Y(n_2815_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2816 (.A1(n_2505_o_0),
    .A2(n_2498_o_0),
    .B(n_2734_o_0),
    .C(n_2591_o_0),
    .D(n_2617_o_0),
    .Y(n_2816_o_0));
 OAI21xp33_ASAP7_75t_R n_2817 (.A1(n_2527_o_0),
    .A2(n_2816_o_0),
    .B(n_2532_o_0),
    .Y(n_2817_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2818 (.A1(n_2815_o_0),
    .A2(n_2527_o_0),
    .B(n_2817_o_0),
    .C(n_2384_o_0),
    .Y(n_2818_o_0));
 AOI21xp33_ASAP7_75t_R n_2819 (.A1(n_2812_o_0),
    .A2(n_2742_o_0),
    .B(n_2818_o_0),
    .Y(n_2819_o_0));
 AOI211xp5_ASAP7_75t_R n_2820 (.A1(n_2810_o_0),
    .A2(n_2385_o_0),
    .B(n_2819_o_0),
    .C(n_2372_o_0),
    .Y(n_2820_o_0));
 AOI21xp33_ASAP7_75t_R n_2821 (.A1(n_2372_o_0),
    .A2(n_2798_o_0),
    .B(n_2820_o_0),
    .Y(n_2821_o_0));
 INVx1_ASAP7_75t_R n_2822 (.A(n_2567_o_0),
    .Y(n_2822_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2823 (.A1(n_2822_o_0),
    .A2(n_2568_o_0),
    .B(net52),
    .C(n_2600_o_0),
    .Y(n_2823_o_0));
 NAND2xp33_ASAP7_75t_R n_2824 (.A(n_2437_o_0),
    .B(n_2459_o_0),
    .Y(n_2824_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2825 (.A1(net75),
    .A2(n_2459_o_0),
    .B(n_2824_o_0),
    .C(n_2507_o_0),
    .Y(n_2825_o_0));
 INVx1_ASAP7_75t_R n_2826 (.A(n_2825_o_0),
    .Y(n_2826_o_0));
 AOI21xp33_ASAP7_75t_R n_2827 (.A1(n_2594_o_0),
    .A2(n_2745_o_0),
    .B(n_2564_o_0),
    .Y(n_2827_o_0));
 AOI21xp33_ASAP7_75t_R n_2828 (.A1(n_2826_o_0),
    .A2(n_2827_o_0),
    .B(n_2384_o_0),
    .Y(n_2828_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2829 (.A1(n_2527_o_0),
    .A2(n_2823_o_0),
    .B(n_2828_o_0),
    .C(n_2532_o_0),
    .Y(n_2829_o_0));
 NOR2xp33_ASAP7_75t_R n_2830 (.A(n_2507_o_0),
    .B(n_2573_o_0),
    .Y(n_2830_o_0));
 OAI22xp33_ASAP7_75t_R n_2831 (.A1(n_2512_o_0),
    .A2(n_2677_o_0),
    .B1(net100),
    .B2(n_2485_o_0),
    .Y(n_2831_o_0));
 AOI21xp33_ASAP7_75t_R n_2832 (.A1(n_2545_o_0),
    .A2(n_2667_o_0),
    .B(n_2527_o_0),
    .Y(n_2832_o_0));
 OAI21xp33_ASAP7_75t_R n_2833 (.A1(n_2415_o_0),
    .A2(net101),
    .B(n_2832_o_0),
    .Y(n_2833_o_0));
 OAI311xp33_ASAP7_75t_R n_2834 (.A1(n_2830_o_0),
    .A2(n_2831_o_0),
    .A3(n_2564_o_0),
    .B1(n_2833_o_0),
    .C1(n_2384_o_0),
    .Y(n_2834_o_0));
 OAI211xp5_ASAP7_75t_R n_2835 (.A1(ld),
    .A2(n_2546_o_0),
    .B(n_2633_o_0),
    .C(n_2415_o_0),
    .Y(n_2835_o_0));
 NAND2xp33_ASAP7_75t_R n_2836 (.A(n_2505_o_0),
    .B(n_2492_o_0),
    .Y(n_2836_o_0));
 NAND3xp33_ASAP7_75t_R n_2837 (.A(n_2745_o_0),
    .B(n_2836_o_0),
    .C(n_2507_o_0),
    .Y(n_2837_o_0));
 AOI21xp33_ASAP7_75t_R n_2838 (.A1(net100),
    .A2(net102),
    .B(n_2507_o_0),
    .Y(n_2838_o_0));
 AOI211xp5_ASAP7_75t_R n_2839 (.A1(n_2732_o_0),
    .A2(n_2507_o_0),
    .B(n_2527_o_0),
    .C(n_2838_o_0),
    .Y(n_2839_o_0));
 AOI31xp33_ASAP7_75t_R n_2840 (.A1(n_2835_o_0),
    .A2(n_2837_o_0),
    .A3(n_2527_o_0),
    .B(n_2839_o_0),
    .Y(n_2840_o_0));
 OAI21xp33_ASAP7_75t_R n_2841 (.A1(n_2505_o_0),
    .A2(n_2437_o_0),
    .B(n_2492_o_0),
    .Y(n_2841_o_0));
 NAND4xp25_ASAP7_75t_R n_2842 (.A(n_2732_o_0),
    .B(n_2841_o_0),
    .C(n_2564_o_0),
    .D(n_2415_o_0),
    .Y(n_2842_o_0));
 AOI21xp33_ASAP7_75t_R n_2843 (.A1(net21),
    .A2(n_2506_o_0),
    .B(n_2507_o_0),
    .Y(n_2843_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2844 (.A1(n_2657_o_0),
    .A2(n_2507_o_0),
    .B(n_2843_o_0),
    .C(n_2527_o_0),
    .Y(n_2844_o_0));
 NAND4xp25_ASAP7_75t_R n_2845 (.A(n_2842_o_0),
    .B(n_2844_o_0),
    .C(n_2609_o_0),
    .D(n_2384_o_0),
    .Y(n_2845_o_0));
 OAI21xp33_ASAP7_75t_R n_2846 (.A1(n_2384_o_0),
    .A2(n_2840_o_0),
    .B(n_2845_o_0),
    .Y(n_2846_o_0));
 AOI221xp5_ASAP7_75t_R n_2847 (.A1(n_2829_o_0),
    .A2(n_2834_o_0),
    .B1(n_2532_o_0),
    .B2(n_2846_o_0),
    .C(n_2372_o_0),
    .Y(n_2847_o_0));
 INVx1_ASAP7_75t_R n_2848 (.A(n_2847_o_0),
    .Y(n_2848_o_0));
 AND2x2_ASAP7_75t_R n_2849 (.A(n_2575_o_0),
    .B(n_2680_o_0),
    .Y(n_2849_o_0));
 NOR2xp33_ASAP7_75t_R n_2850 (.A(n_2668_o_0),
    .B(n_2675_o_0),
    .Y(n_2850_o_0));
 OAI221xp5_ASAP7_75t_R n_2851 (.A1(net21),
    .A2(n_2506_o_0),
    .B1(net52),
    .B2(n_2746_o_0),
    .C(n_2527_o_0),
    .Y(n_2851_o_0));
 OAI31xp33_ASAP7_75t_R n_2852 (.A1(n_2527_o_0),
    .A2(n_2849_o_0),
    .A3(n_2850_o_0),
    .B(n_2851_o_0),
    .Y(n_2852_o_0));
 OAI222xp33_ASAP7_75t_R n_2853 (.A1(n_2585_o_0),
    .A2(n_2702_o_0),
    .B1(n_2773_o_0),
    .B2(net21),
    .C1(n_2485_o_0),
    .C2(n_2510_o_0),
    .Y(n_2853_o_0));
 OAI21xp33_ASAP7_75t_R n_2854 (.A1(net21),
    .A2(n_2461_o_0),
    .B(n_2415_o_0),
    .Y(n_2854_o_0));
 AOI31xp33_ASAP7_75t_R n_2855 (.A1(n_2507_o_0),
    .A2(n_2616_o_0),
    .A3(n_2625_o_0),
    .B(n_2527_o_0),
    .Y(n_2855_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2856 (.A1(net21),
    .A2(n_2585_o_0),
    .B(n_2854_o_0),
    .C(n_2855_o_0),
    .Y(n_2856_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2857 (.A1(n_2564_o_0),
    .A2(n_2853_o_0),
    .B(n_2856_o_0),
    .C(n_2384_o_0),
    .Y(n_2857_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2858 (.A1(n_2384_o_0),
    .A2(n_2852_o_0),
    .B(n_2857_o_0),
    .C(n_2532_o_0),
    .Y(n_2858_o_0));
 NAND3xp33_ASAP7_75t_R n_2859 (.A(n_2616_o_0),
    .B(n_2690_o_0),
    .C(n_2507_o_0),
    .Y(n_2859_o_0));
 OAI31xp33_ASAP7_75t_R n_2860 (.A1(n_2507_o_0),
    .A2(n_2782_o_0),
    .A3(n_2645_o_0),
    .B(n_2859_o_0),
    .Y(n_2860_o_0));
 AOI211xp5_ASAP7_75t_R n_2861 (.A1(n_2415_o_0),
    .A2(net102),
    .B(net101),
    .C(n_2505_o_0),
    .Y(n_2861_o_0));
 AOI21xp33_ASAP7_75t_R n_2862 (.A1(n_2507_o_0),
    .A2(n_2661_o_0),
    .B(n_2861_o_0),
    .Y(n_2862_o_0));
 AOI31xp33_ASAP7_75t_R n_2863 (.A1(n_2564_o_0),
    .A2(n_2862_o_0),
    .A3(n_2835_o_0),
    .B(n_2384_o_0),
    .Y(n_2863_o_0));
 OAI21xp33_ASAP7_75t_R n_2864 (.A1(n_2564_o_0),
    .A2(n_2860_o_0),
    .B(n_2863_o_0),
    .Y(n_2864_o_0));
 AOI21xp33_ASAP7_75t_R n_2865 (.A1(net102),
    .A2(net21),
    .B(net100),
    .Y(n_2865_o_0));
 AOI211xp5_ASAP7_75t_R n_2866 (.A1(n_2507_o_0),
    .A2(n_2865_o_0),
    .B(n_2825_o_0),
    .C(n_2564_o_0),
    .Y(n_2866_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2867 (.A1(n_2666_o_0),
    .A2(n_2675_o_0),
    .B(n_2764_o_0),
    .C(n_2527_o_0),
    .Y(n_2867_o_0));
 OAI21xp33_ASAP7_75t_R n_2868 (.A1(n_2866_o_0),
    .A2(n_2867_o_0),
    .B(n_2384_o_0),
    .Y(n_2868_o_0));
 NAND3xp33_ASAP7_75t_R n_2869 (.A(n_2864_o_0),
    .B(n_2396_o_0),
    .C(n_2868_o_0),
    .Y(n_2869_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2870 (.A1(n_2858_o_0),
    .A2(n_2869_o_0),
    .B(n_2847_o_0),
    .C(n_2372_o_0),
    .Y(n_2870_o_0));
 OAI21xp33_ASAP7_75t_R n_2871 (.A1(n_2372_o_0),
    .A2(n_2848_o_0),
    .B(n_2870_o_0),
    .Y(n_2871_o_0));
 OAI211xp5_ASAP7_75t_R n_2872 (.A1(net52),
    .A2(net100),
    .B(n_2826_o_0),
    .C(n_2532_o_0),
    .Y(n_2872_o_0));
 NAND2xp33_ASAP7_75t_R n_2873 (.A(n_2741_o_0),
    .B(n_2396_o_0),
    .Y(n_2873_o_0));
 AO21x1_ASAP7_75t_R n_2874 (.A1(n_2544_o_0),
    .A2(n_2598_o_0),
    .B(n_2873_o_0),
    .Y(n_2874_o_0));
 AOI21xp33_ASAP7_75t_R n_2875 (.A1(n_2872_o_0),
    .A2(n_2874_o_0),
    .B(n_2527_o_0),
    .Y(n_2875_o_0));
 AOI21xp33_ASAP7_75t_R n_2876 (.A1(net101),
    .A2(n_2460_o_0),
    .B(n_2415_o_0),
    .Y(n_2876_o_0));
 AOI22xp33_ASAP7_75t_R n_2877 (.A1(n_2774_o_0),
    .A2(n_2876_o_0),
    .B1(n_2584_o_0),
    .B2(n_2514_o_0),
    .Y(n_2877_o_0));
 OAI21xp33_ASAP7_75t_R n_2878 (.A1(n_2585_o_0),
    .A2(n_2702_o_0),
    .B(n_2396_o_0),
    .Y(n_2878_o_0));
 AO21x1_ASAP7_75t_R n_2879 (.A1(n_2734_o_0),
    .A2(n_2562_o_0),
    .B(n_2878_o_0),
    .Y(n_2879_o_0));
 OAI21xp33_ASAP7_75t_R n_2880 (.A1(n_2396_o_0),
    .A2(n_2877_o_0),
    .B(n_2879_o_0),
    .Y(n_2880_o_0));
 OAI21xp33_ASAP7_75t_R n_2881 (.A1(n_2564_o_0),
    .A2(n_2880_o_0),
    .B(n_2385_o_0),
    .Y(n_2881_o_0));
 NAND3xp33_ASAP7_75t_R n_2882 (.A(n_2616_o_0),
    .B(net52),
    .C(n_2625_o_0),
    .Y(n_2882_o_0));
 AOI21xp33_ASAP7_75t_R n_2883 (.A1(n_2594_o_0),
    .A2(n_2710_o_0),
    .B(n_2564_o_0),
    .Y(n_2883_o_0));
 AO21x1_ASAP7_75t_R n_2884 (.A1(n_2882_o_0),
    .A2(n_2883_o_0),
    .B(n_2396_o_0),
    .Y(n_2884_o_0));
 NOR2xp33_ASAP7_75t_R n_2885 (.A(n_2512_o_0),
    .B(n_2813_o_0),
    .Y(n_2885_o_0));
 NOR4xp25_ASAP7_75t_R n_2886 (.A(n_2885_o_0),
    .B(n_2583_o_0),
    .C(n_2508_o_0),
    .D(n_2527_o_0),
    .Y(n_2886_o_0));
 INVx1_ASAP7_75t_R n_2887 (.A(n_2841_o_0),
    .Y(n_2887_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2888 (.A1(n_2507_o_0),
    .A2(n_2511_o_0),
    .B(n_2887_o_0),
    .C(n_2527_o_0),
    .Y(n_2888_o_0));
 AOI21xp33_ASAP7_75t_R n_2889 (.A1(n_2415_o_0),
    .A2(n_2662_o_0),
    .B(n_2527_o_0),
    .Y(n_2889_o_0));
 OAI321xp33_ASAP7_75t_R n_2890 (.A1(net52),
    .A2(net21),
    .A3(n_2773_o_0),
    .B1(n_2702_o_0),
    .B2(net102),
    .C(n_2889_o_0),
    .Y(n_2890_o_0));
 AOI31xp33_ASAP7_75t_R n_2891 (.A1(n_2888_o_0),
    .A2(n_2890_o_0),
    .A3(n_2396_o_0),
    .B(n_2385_o_0),
    .Y(n_2891_o_0));
 OAI21xp33_ASAP7_75t_R n_2892 (.A1(n_2884_o_0),
    .A2(n_2886_o_0),
    .B(n_2891_o_0),
    .Y(n_2892_o_0));
 OAI21xp33_ASAP7_75t_R n_2893 (.A1(n_2875_o_0),
    .A2(n_2881_o_0),
    .B(n_2892_o_0),
    .Y(n_2893_o_0));
 NAND3xp33_ASAP7_75t_R n_2894 (.A(n_2543_o_0),
    .B(n_2686_o_0),
    .C(n_2507_o_0),
    .Y(n_2894_o_0));
 OAI31xp33_ASAP7_75t_R n_2895 (.A1(n_2507_o_0),
    .A2(n_2782_o_0),
    .A3(n_2699_o_0),
    .B(n_2894_o_0),
    .Y(n_2895_o_0));
 AOI21xp33_ASAP7_75t_R n_2896 (.A1(n_2396_o_0),
    .A2(n_2895_o_0),
    .B(n_2564_o_0),
    .Y(n_2896_o_0));
 OAI22xp33_ASAP7_75t_R n_2897 (.A1(n_2813_o_0),
    .A2(net52),
    .B1(n_2510_o_0),
    .B2(n_2485_o_0),
    .Y(n_2897_o_0));
 NAND2xp33_ASAP7_75t_R n_2898 (.A(n_2532_o_0),
    .B(n_2897_o_0),
    .Y(n_2898_o_0));
 AO21x1_ASAP7_75t_R n_2899 (.A1(n_2507_o_0),
    .A2(n_2773_o_0),
    .B(n_2685_o_0),
    .Y(n_2899_o_0));
 AOI31xp33_ASAP7_75t_R n_2900 (.A1(n_2415_o_0),
    .A2(n_2510_o_0),
    .A3(net21),
    .B(n_2653_o_0),
    .Y(n_2900_o_0));
 NAND3xp33_ASAP7_75t_R n_2901 (.A(n_2900_o_0),
    .B(n_2806_o_0),
    .C(n_2532_o_0),
    .Y(n_2901_o_0));
 OAI21xp33_ASAP7_75t_R n_2902 (.A1(n_2532_o_0),
    .A2(n_2899_o_0),
    .B(n_2901_o_0),
    .Y(n_2902_o_0));
 AOI22xp33_ASAP7_75t_R n_2903 (.A1(n_2896_o_0),
    .A2(n_2898_o_0),
    .B1(n_2564_o_0),
    .B2(n_2902_o_0),
    .Y(n_2903_o_0));
 AOI31xp33_ASAP7_75t_R n_2904 (.A1(n_2507_o_0),
    .A2(n_2548_o_0),
    .A3(n_2543_o_0),
    .B(n_2396_o_0),
    .Y(n_2904_o_0));
 OAI21xp33_ASAP7_75t_R n_2905 (.A1(n_2554_o_0),
    .A2(n_2746_o_0),
    .B(n_2904_o_0),
    .Y(n_2905_o_0));
 AOI21xp33_ASAP7_75t_R n_2906 (.A1(n_2545_o_0),
    .A2(n_2685_o_0),
    .B(n_2532_o_0),
    .Y(n_2906_o_0));
 OAI31xp33_ASAP7_75t_R n_2907 (.A1(net52),
    .A2(net101),
    .A3(n_2576_o_0),
    .B(n_2906_o_0),
    .Y(n_2907_o_0));
 NAND3xp33_ASAP7_75t_R n_2908 (.A(n_2905_o_0),
    .B(n_2907_o_0),
    .C(n_2527_o_0),
    .Y(n_2908_o_0));
 AOI22xp33_ASAP7_75t_R n_2909 (.A1(n_2710_o_0),
    .A2(n_2680_o_0),
    .B1(net102),
    .B2(n_2793_o_0),
    .Y(n_2909_o_0));
 OAI21xp33_ASAP7_75t_R n_2910 (.A1(net52),
    .A2(n_2632_o_0),
    .B(n_2909_o_0),
    .Y(n_2910_o_0));
 AOI21xp33_ASAP7_75t_R n_2911 (.A1(n_2568_o_0),
    .A2(n_2667_o_0),
    .B(n_2396_o_0),
    .Y(n_2911_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2912 (.A1(net52),
    .A2(n_2498_o_0),
    .B(n_2911_o_0),
    .C(n_2527_o_0),
    .Y(n_2912_o_0));
 OAI21xp33_ASAP7_75t_R n_2913 (.A1(n_2910_o_0),
    .A2(n_2532_o_0),
    .B(n_2912_o_0),
    .Y(n_2913_o_0));
 AOI31xp33_ASAP7_75t_R n_2914 (.A1(n_2384_o_0),
    .A2(n_2908_o_0),
    .A3(n_2913_o_0),
    .B(n_2372_o_0),
    .Y(n_2914_o_0));
 OAI21xp33_ASAP7_75t_R n_2915 (.A1(n_2903_o_0),
    .A2(n_2384_o_0),
    .B(n_2914_o_0),
    .Y(n_2915_o_0));
 OAI21xp33_ASAP7_75t_R n_2916 (.A1(n_2373_o_0),
    .A2(n_2893_o_0),
    .B(n_2915_o_0),
    .Y(n_2916_o_0));
 INVx1_ASAP7_75t_R n_2917 (.A(n_2623_o_0),
    .Y(n_2917_o_0));
 AOI21xp33_ASAP7_75t_R n_2918 (.A1(n_2917_o_0),
    .A2(n_2837_o_0),
    .B(n_2564_o_0),
    .Y(n_2918_o_0));
 OR3x1_ASAP7_75t_R n_2919 (.A(n_2918_o_0),
    .B(n_2736_o_0),
    .C(n_2532_o_0),
    .Y(n_2919_o_0));
 AOI21xp33_ASAP7_75t_R n_2920 (.A1(net100),
    .A2(net101),
    .B(n_2677_o_0),
    .Y(n_2920_o_0));
 INVx1_ASAP7_75t_R n_2921 (.A(n_2554_o_0),
    .Y(n_2921_o_0));
 AOI22xp33_ASAP7_75t_R n_2922 (.A1(n_2920_o_0),
    .A2(n_2507_o_0),
    .B1(n_2921_o_0),
    .B2(n_2745_o_0),
    .Y(n_2922_o_0));
 AOI31xp33_ASAP7_75t_R n_2923 (.A1(n_2507_o_0),
    .A2(n_2561_o_0),
    .A3(n_2543_o_0),
    .B(n_2564_o_0),
    .Y(n_2923_o_0));
 AOI21xp33_ASAP7_75t_R n_2924 (.A1(n_2613_o_0),
    .A2(n_2923_o_0),
    .B(n_2396_o_0),
    .Y(n_2924_o_0));
 OAI21xp33_ASAP7_75t_R n_2925 (.A1(n_2527_o_0),
    .A2(n_2922_o_0),
    .B(n_2924_o_0),
    .Y(n_2925_o_0));
 OAI311xp33_ASAP7_75t_R n_2926 (.A1(net21),
    .A2(n_2540_o_0),
    .A3(n_2538_o_0),
    .B1(n_2598_o_0),
    .C1(n_2415_o_0),
    .Y(n_2926_o_0));
 OAI31xp33_ASAP7_75t_R n_2927 (.A1(n_2593_o_0),
    .A2(n_2555_o_0),
    .A3(net52),
    .B(n_2926_o_0),
    .Y(n_2927_o_0));
 OAI21xp33_ASAP7_75t_R n_2928 (.A1(n_2507_o_0),
    .A2(n_2662_o_0),
    .B(n_2527_o_0),
    .Y(n_2928_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2929 (.A1(n_2927_o_0),
    .A2(n_2564_o_0),
    .B(n_2396_o_0),
    .C(n_2928_o_0),
    .Y(n_2929_o_0));
 OAI221xp5_ASAP7_75t_R n_2930 (.A1(n_2507_o_0),
    .A2(n_2662_o_0),
    .B1(n_2396_o_0),
    .B2(n_2716_o_0),
    .C(n_2527_o_0),
    .Y(n_2930_o_0));
 AOI31xp33_ASAP7_75t_R n_2931 (.A1(n_2507_o_0),
    .A2(n_2616_o_0),
    .A3(n_2674_o_0),
    .B(n_2564_o_0),
    .Y(n_2931_o_0));
 OAI21xp33_ASAP7_75t_R n_2932 (.A1(n_2774_o_0),
    .A2(n_2507_o_0),
    .B(n_2931_o_0),
    .Y(n_2932_o_0));
 AOI31xp33_ASAP7_75t_R n_2933 (.A1(n_2642_o_0),
    .A2(n_2616_o_0),
    .A3(n_2507_o_0),
    .B(n_2527_o_0),
    .Y(n_2933_o_0));
 OAI21xp33_ASAP7_75t_R n_2934 (.A1(n_2666_o_0),
    .A2(n_2743_o_0),
    .B(n_2933_o_0),
    .Y(n_2934_o_0));
 AOI21xp33_ASAP7_75t_R n_2935 (.A1(n_2932_o_0),
    .A2(n_2934_o_0),
    .B(n_2532_o_0),
    .Y(n_2935_o_0));
 AOI211xp5_ASAP7_75t_R n_2936 (.A1(n_2929_o_0),
    .A2(n_2930_o_0),
    .B(n_2935_o_0),
    .C(n_2373_o_0),
    .Y(n_2936_o_0));
 AOI31xp33_ASAP7_75t_R n_2937 (.A1(n_2373_o_0),
    .A2(n_2919_o_0),
    .A3(n_2925_o_0),
    .B(n_2936_o_0),
    .Y(n_2937_o_0));
 INVx1_ASAP7_75t_R n_2938 (.A(n_2814_o_0),
    .Y(n_2938_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2939 (.A1(net52),
    .A2(n_2699_o_0),
    .B(n_2938_o_0),
    .C(n_2564_o_0),
    .Y(n_2939_o_0));
 OAI21xp33_ASAP7_75t_R n_2940 (.A1(net52),
    .A2(n_2637_o_0),
    .B(n_2549_o_0),
    .Y(n_2940_o_0));
 AOI21xp33_ASAP7_75t_R n_2941 (.A1(n_2527_o_0),
    .A2(n_2940_o_0),
    .B(n_2532_o_0),
    .Y(n_2941_o_0));
 NAND3xp33_ASAP7_75t_R n_2942 (.A(n_2695_o_0),
    .B(n_2591_o_0),
    .C(n_2507_o_0),
    .Y(n_2942_o_0));
 AOI21xp33_ASAP7_75t_R n_2943 (.A1(n_2710_o_0),
    .A2(n_2921_o_0),
    .B(n_2527_o_0),
    .Y(n_2943_o_0));
 AOI21xp33_ASAP7_75t_R n_2944 (.A1(n_2507_o_0),
    .A2(n_2568_o_0),
    .B(n_2698_o_0),
    .Y(n_2944_o_0));
 NOR3xp33_ASAP7_75t_R n_2945 (.A(n_2944_o_0),
    .B(n_2564_o_0),
    .C(n_2643_o_0),
    .Y(n_2945_o_0));
 AOI211xp5_ASAP7_75t_R n_2946 (.A1(n_2942_o_0),
    .A2(n_2943_o_0),
    .B(n_2945_o_0),
    .C(n_2396_o_0),
    .Y(n_2946_o_0));
 AOI21xp33_ASAP7_75t_R n_2947 (.A1(n_2939_o_0),
    .A2(n_2941_o_0),
    .B(n_2946_o_0),
    .Y(n_2947_o_0));
 AOI22xp33_ASAP7_75t_R n_2948 (.A1(n_2793_o_0),
    .A2(n_2574_o_0),
    .B1(n_2804_o_0),
    .B2(n_2576_o_0),
    .Y(n_2948_o_0));
 OAI21xp33_ASAP7_75t_R n_2949 (.A1(n_2507_o_0),
    .A2(n_2573_o_0),
    .B(n_2948_o_0),
    .Y(n_2949_o_0));
 AOI21xp33_ASAP7_75t_R n_2950 (.A1(n_2584_o_0),
    .A2(n_2836_o_0),
    .B(net52),
    .Y(n_2950_o_0));
 OAI21xp33_ASAP7_75t_R n_2951 (.A1(n_2507_o_0),
    .A2(net100),
    .B(n_2564_o_0),
    .Y(n_2951_o_0));
 OAI22xp33_ASAP7_75t_R n_2952 (.A1(n_2949_o_0),
    .A2(n_2564_o_0),
    .B1(n_2950_o_0),
    .B2(n_2951_o_0),
    .Y(n_2952_o_0));
 OAI211xp5_ASAP7_75t_R n_2953 (.A1(net21),
    .A2(n_2574_o_0),
    .B(n_2657_o_0),
    .C(n_2507_o_0),
    .Y(n_2953_o_0));
 AOI21xp33_ASAP7_75t_R n_2954 (.A1(n_2745_o_0),
    .A2(n_2698_o_0),
    .B(n_2527_o_0),
    .Y(n_2954_o_0));
 AOI21xp33_ASAP7_75t_R n_2955 (.A1(n_2953_o_0),
    .A2(n_2954_o_0),
    .B(n_2532_o_0),
    .Y(n_2955_o_0));
 INVx1_ASAP7_75t_R n_2956 (.A(n_2566_o_0),
    .Y(n_2956_o_0));
 OAI31xp33_ASAP7_75t_R n_2957 (.A1(n_2415_o_0),
    .A2(n_2773_o_0),
    .A3(net21),
    .B(n_2527_o_0),
    .Y(n_2957_o_0));
 AOI21xp33_ASAP7_75t_R n_2958 (.A1(n_2956_o_0),
    .A2(n_2732_o_0),
    .B(n_2957_o_0),
    .Y(n_2958_o_0));
 OAI21xp33_ASAP7_75t_R n_2959 (.A1(net102),
    .A2(n_2702_o_0),
    .B(n_2958_o_0),
    .Y(n_2959_o_0));
 AOI21xp33_ASAP7_75t_R n_2960 (.A1(n_2955_o_0),
    .A2(n_2959_o_0),
    .B(n_2373_o_0),
    .Y(n_2960_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2961 (.A1(n_2952_o_0),
    .A2(n_2396_o_0),
    .B(n_2960_o_0),
    .C(n_2385_o_0),
    .Y(n_2961_o_0));
 OAI21xp33_ASAP7_75t_R n_2962 (.A1(n_2947_o_0),
    .A2(n_2372_o_0),
    .B(n_2961_o_0),
    .Y(n_2962_o_0));
 OAI21xp33_ASAP7_75t_R n_2963 (.A1(n_2384_o_0),
    .A2(n_2937_o_0),
    .B(n_2962_o_0),
    .Y(n_2963_o_0));
 OAI21xp33_ASAP7_75t_R n_2964 (.A1(n_2789_o_0),
    .A2(n_2592_o_0),
    .B(n_2807_o_0),
    .Y(n_2964_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_2965 (.A1(n_2668_o_0),
    .A2(n_2691_o_0),
    .B(n_2954_o_0),
    .C(n_2532_o_0),
    .Y(n_2965_o_0));
 OA21x2_ASAP7_75t_R n_2966 (.A1(n_2964_o_0),
    .A2(n_2564_o_0),
    .B(n_2965_o_0),
    .Y(n_2966_o_0));
 AND3x1_ASAP7_75t_R n_2967 (.A(n_2837_o_0),
    .B(n_2854_o_0),
    .C(n_2564_o_0),
    .Y(n_2967_o_0));
 OA211x2_ASAP7_75t_R n_2968 (.A1(net21),
    .A2(n_2506_o_0),
    .B(n_2657_o_0),
    .C(n_2507_o_0),
    .Y(n_2968_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_2969 (.A1(n_2514_o_0),
    .A2(n_2616_o_0),
    .B(n_2968_o_0),
    .C(n_2532_o_0),
    .D(n_2564_o_0),
    .Y(n_2969_o_0));
 NOR2xp33_ASAP7_75t_R n_2970 (.A(n_2527_o_0),
    .B(n_2532_o_0),
    .Y(n_2970_o_0));
 OAI31xp33_ASAP7_75t_R n_2971 (.A1(n_2967_o_0),
    .A2(n_2969_o_0),
    .A3(n_2970_o_0),
    .B(n_2384_o_0),
    .Y(n_2971_o_0));
 INVx1_ASAP7_75t_R n_2972 (.A(n_2876_o_0),
    .Y(n_2972_o_0));
 AOI22xp33_ASAP7_75t_R n_2973 (.A1(n_2783_o_0),
    .A2(n_2657_o_0),
    .B1(n_2616_o_0),
    .B2(n_2507_o_0),
    .Y(n_2973_o_0));
 OAI21xp33_ASAP7_75t_R n_2974 (.A1(n_2564_o_0),
    .A2(n_2973_o_0),
    .B(n_2396_o_0),
    .Y(n_2974_o_0));
 AOI21xp33_ASAP7_75t_R n_2975 (.A1(n_2972_o_0),
    .A2(n_2889_o_0),
    .B(n_2974_o_0),
    .Y(n_2975_o_0));
 NAND2xp33_ASAP7_75t_R n_2976 (.A(n_2657_o_0),
    .B(n_2921_o_0),
    .Y(n_2976_o_0));
 OAI31xp33_ASAP7_75t_R n_2977 (.A1(n_2569_o_0),
    .A2(n_2718_o_0),
    .A3(net52),
    .B(n_2976_o_0),
    .Y(n_2977_o_0));
 OAI21xp33_ASAP7_75t_R n_2978 (.A1(net102),
    .A2(n_2507_o_0),
    .B(n_2527_o_0),
    .Y(n_2978_o_0));
 OAI21xp33_ASAP7_75t_R n_2979 (.A1(n_2978_o_0),
    .A2(n_2850_o_0),
    .B(n_2532_o_0),
    .Y(n_2979_o_0));
 AOI21xp33_ASAP7_75t_R n_2980 (.A1(n_2564_o_0),
    .A2(n_2977_o_0),
    .B(n_2979_o_0),
    .Y(n_2980_o_0));
 OAI21xp33_ASAP7_75t_R n_2981 (.A1(n_2975_o_0),
    .A2(n_2980_o_0),
    .B(n_2385_o_0),
    .Y(n_2981_o_0));
 OAI21xp33_ASAP7_75t_R n_2982 (.A1(n_2966_o_0),
    .A2(n_2971_o_0),
    .B(n_2981_o_0),
    .Y(n_2982_o_0));
 OAI211xp5_ASAP7_75t_R n_2983 (.A1(n_2585_o_0),
    .A2(net101),
    .B(n_2543_o_0),
    .C(n_2507_o_0),
    .Y(n_2983_o_0));
 OAI31xp33_ASAP7_75t_R n_2984 (.A1(n_2507_o_0),
    .A2(n_2619_o_0),
    .A3(n_2643_o_0),
    .B(n_2983_o_0),
    .Y(n_2984_o_0));
 AOI211xp5_ASAP7_75t_R n_2985 (.A1(net52),
    .A2(n_2635_o_0),
    .B(n_2831_o_0),
    .C(n_2396_o_0),
    .Y(n_2985_o_0));
 AOI21xp33_ASAP7_75t_R n_2986 (.A1(n_2396_o_0),
    .A2(n_2984_o_0),
    .B(n_2985_o_0),
    .Y(n_2986_o_0));
 OAI21xp33_ASAP7_75t_R n_2987 (.A1(net52),
    .A2(n_2684_o_0),
    .B(n_2606_o_0),
    .Y(n_2987_o_0));
 AOI211xp5_ASAP7_75t_R n_2988 (.A1(net52),
    .A2(n_2592_o_0),
    .B(n_2987_o_0),
    .C(n_2532_o_0),
    .Y(n_2988_o_0));
 NOR3xp33_ASAP7_75t_R n_2989 (.A(n_2506_o_0),
    .B(n_2507_o_0),
    .C(n_2492_o_0),
    .Y(n_2989_o_0));
 AOI211xp5_ASAP7_75t_R n_2990 (.A1(n_2507_o_0),
    .A2(n_2460_o_0),
    .B(n_2989_o_0),
    .C(n_2396_o_0),
    .Y(n_2990_o_0));
 OAI31xp33_ASAP7_75t_R n_2991 (.A1(n_2527_o_0),
    .A2(n_2988_o_0),
    .A3(n_2990_o_0),
    .B(n_2385_o_0),
    .Y(n_2991_o_0));
 OA21x2_ASAP7_75t_R n_2992 (.A1(net21),
    .A2(n_2506_o_0),
    .B(n_2657_o_0),
    .Y(n_2992_o_0));
 NAND2xp33_ASAP7_75t_R n_2993 (.A(net21),
    .B(n_2773_o_0),
    .Y(n_2993_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2994 (.A1(n_2993_o_0),
    .A2(n_2543_o_0),
    .B(net52),
    .C(n_2564_o_0),
    .Y(n_2994_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2995 (.A1(n_2461_o_0),
    .A2(net21),
    .B(n_2735_o_0),
    .C(n_2827_o_0),
    .Y(n_2995_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_2996 (.A1(n_2992_o_0),
    .A2(net52),
    .B(n_2994_o_0),
    .C(n_2995_o_0),
    .Y(n_2996_o_0));
 OAI21xp33_ASAP7_75t_R n_2997 (.A1(n_2510_o_0),
    .A2(n_2507_o_0),
    .B(n_2527_o_0),
    .Y(n_2997_o_0));
 AOI21xp33_ASAP7_75t_R n_2998 (.A1(n_2505_o_0),
    .A2(n_2793_o_0),
    .B(n_2989_o_0),
    .Y(n_2998_o_0));
 AOI31xp33_ASAP7_75t_R n_2999 (.A1(n_2564_o_0),
    .A2(n_2573_o_0),
    .A3(n_2998_o_0),
    .B(n_2532_o_0),
    .Y(n_2999_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3000 (.A1(n_2950_o_0),
    .A2(n_2997_o_0),
    .B(n_2999_o_0),
    .C(n_2385_o_0),
    .Y(n_3000_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3001 (.A1(n_2396_o_0),
    .A2(n_2996_o_0),
    .B(n_3000_o_0),
    .C(n_2373_o_0),
    .Y(n_3001_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3002 (.A1(n_2527_o_0),
    .A2(n_2986_o_0),
    .B(n_2991_o_0),
    .C(n_3001_o_0),
    .Y(n_3002_o_0));
 OAI21xp33_ASAP7_75t_R n_3003 (.A1(n_2372_o_0),
    .A2(n_2982_o_0),
    .B(n_3002_o_0),
    .Y(n_3003_o_0));
 XNOR2xp5_ASAP7_75t_R n_3004 (.A(_01000_),
    .B(_01040_),
    .Y(n_3004_o_0));
 XNOR2xp5_ASAP7_75t_R n_3005 (.A(_01081_),
    .B(_01120_),
    .Y(n_3005_o_0));
 XNOR2xp5_ASAP7_75t_R n_3006 (.A(_01041_),
    .B(n_3005_o_0),
    .Y(n_3006_o_0));
 XOR2xp5_ASAP7_75t_R n_3007 (.A(n_3004_o_0),
    .B(n_3006_o_0),
    .Y(n_3007_o_0));
 NOR2xp33_ASAP7_75t_R n_3008 (.A(_00651_),
    .B(net),
    .Y(n_3008_o_0));
 AOI21xp33_ASAP7_75t_R n_3009 (.A1(net39),
    .A2(n_3007_o_0),
    .B(n_3008_o_0),
    .Y(n_3009_o_0));
 XNOR2xp5_ASAP7_75t_R n_3010 (.A(_00889_),
    .B(n_3009_o_0),
    .Y(n_3010_o_0));
 XOR2xp5_ASAP7_75t_R n_3011 (.A(_01002_),
    .B(_01042_),
    .Y(n_3011_o_0));
 XNOR2xp5_ASAP7_75t_R n_3012 (.A(_00642_),
    .B(_00643_),
    .Y(n_3012_o_0));
 XNOR2xp5_ASAP7_75t_R n_3013 (.A(_01043_),
    .B(n_3012_o_0),
    .Y(n_3013_o_0));
 NAND2xp33_ASAP7_75t_R n_3014 (.A(n_3011_o_0),
    .B(n_3013_o_0),
    .Y(n_3014_o_0));
 OAI21xp33_ASAP7_75t_R n_3015 (.A1(n_3011_o_0),
    .A2(n_3013_o_0),
    .B(n_3014_o_0),
    .Y(n_3015_o_0));
 NOR2xp33_ASAP7_75t_R n_3016 (.A(_00649_),
    .B(net),
    .Y(n_3016_o_0));
 AOI211xp5_ASAP7_75t_R n_3017 (.A1(n_3015_o_0),
    .A2(net),
    .B(_00891_),
    .C(n_3016_o_0),
    .Y(n_3017_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3018 (.A1(n_3015_o_0),
    .A2(net),
    .B(n_3016_o_0),
    .C(_00891_),
    .Y(n_3018_o_0));
 INVx1_ASAP7_75t_R n_3019 (.A(n_3018_o_0),
    .Y(n_3019_o_0));
 NOR2xp33_ASAP7_75t_R n_3020 (.A(n_3017_o_0),
    .B(n_3019_o_0),
    .Y(n_3020_o_0));
 INVx3_ASAP7_75t_R n_3021 (.A(_00858_),
    .Y(n_3021_o_0));
 XNOR2xp5_ASAP7_75t_R n_3022 (.A(_00998_),
    .B(_01003_),
    .Y(n_3022_o_0));
 NAND2xp33_ASAP7_75t_R n_3023 (.A(_01039_),
    .B(n_3022_o_0),
    .Y(n_3023_o_0));
 OAI21xp33_ASAP7_75t_R n_3024 (.A1(_01039_),
    .A2(n_3022_o_0),
    .B(n_3023_o_0),
    .Y(n_3024_o_0));
 XNOR2xp5_ASAP7_75t_R n_3025 (.A(_01038_),
    .B(_01043_),
    .Y(n_3025_o_0));
 XNOR2xp5_ASAP7_75t_R n_3026 (.A(_01079_),
    .B(_01118_),
    .Y(n_3026_o_0));
 XNOR2xp5_ASAP7_75t_R n_3027 (.A(n_3025_o_0),
    .B(n_3026_o_0),
    .Y(n_3027_o_0));
 XNOR2xp5_ASAP7_75t_R n_3028 (.A(n_3024_o_0),
    .B(n_3027_o_0),
    .Y(n_3028_o_0));
 NOR2xp33_ASAP7_75t_R n_3029 (.A(_00653_),
    .B(_00858_),
    .Y(n_3029_o_0));
 INVx1_ASAP7_75t_R n_3030 (.A(n_3029_o_0),
    .Y(n_3030_o_0));
 OAI21xp33_ASAP7_75t_R n_3031 (.A1(net3),
    .A2(n_3028_o_0),
    .B(n_3030_o_0),
    .Y(n_3031_o_0));
 XOR2xp5_ASAP7_75t_R n_3032 (.A(n_3024_o_0),
    .B(n_3027_o_0),
    .Y(n_3032_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3033 (.A1(n_3032_o_0),
    .A2(net),
    .B(n_3029_o_0),
    .C(_00887_),
    .Y(n_3033_o_0));
 OAI21xp5_ASAP7_75t_R n_3034 (.A1(_00887_),
    .A2(n_3031_o_0),
    .B(n_3033_o_0),
    .Y(n_3034_o_0));
 XNOR2xp5_ASAP7_75t_R n_3035 (.A(_00997_),
    .B(_01037_),
    .Y(n_3035_o_0));
 INVx1_ASAP7_75t_R n_3036 (.A(n_3035_o_0),
    .Y(n_3036_o_0));
 XNOR2xp5_ASAP7_75t_R n_3037 (.A(_01078_),
    .B(_01117_),
    .Y(n_3037_o_0));
 XNOR2xp5_ASAP7_75t_R n_3038 (.A(_01038_),
    .B(n_3037_o_0),
    .Y(n_3038_o_0));
 OAI21xp33_ASAP7_75t_R n_3039 (.A1(n_3036_o_0),
    .A2(n_3038_o_0),
    .B(net39),
    .Y(n_3039_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3040 (.A1(n_3036_o_0),
    .A2(n_3038_o_0),
    .B(n_3039_o_0),
    .C(_00886_),
    .Y(n_3040_o_0));
 XNOR2xp5_ASAP7_75t_R n_3041 (.A(n_3035_o_0),
    .B(n_3038_o_0),
    .Y(n_3041_o_0));
 OAI21xp33_ASAP7_75t_R n_3042 (.A1(_00492_),
    .A2(net39),
    .B(n_2464_o_0),
    .Y(n_3042_o_0));
 INVx1_ASAP7_75t_R n_3043 (.A(n_3042_o_0),
    .Y(n_3043_o_0));
 OAI21xp33_ASAP7_75t_R n_3044 (.A1(n_3021_o_0),
    .A2(n_3041_o_0),
    .B(n_3043_o_0),
    .Y(n_3044_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3045 (.A1(net3),
    .A2(_00492_),
    .B(n_3040_o_0),
    .C(n_3044_o_0),
    .Y(n_3045_o_0));
 XNOR2xp5_ASAP7_75t_R n_3046 (.A(_01036_),
    .B(_01076_),
    .Y(n_3046_o_0));
 INVx1_ASAP7_75t_R n_3047 (.A(n_3046_o_0),
    .Y(n_3047_o_0));
 XNOR2xp5_ASAP7_75t_R n_3048 (.A(_01003_),
    .B(_01043_),
    .Y(n_3048_o_0));
 XNOR2xp5_ASAP7_75t_R n_3049 (.A(_01115_),
    .B(n_3048_o_0),
    .Y(n_3049_o_0));
 INVx1_ASAP7_75t_R n_3050 (.A(_01115_),
    .Y(n_3050_o_0));
 NAND2xp33_ASAP7_75t_R n_3051 (.A(n_3050_o_0),
    .B(n_3048_o_0),
    .Y(n_3051_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3052 (.A1(n_3048_o_0),
    .A2(n_3050_o_0),
    .B(n_3051_o_0),
    .C(n_3047_o_0),
    .Y(n_3052_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3053 (.A1(n_3047_o_0),
    .A2(n_3049_o_0),
    .B(n_3052_o_0),
    .C(net39),
    .Y(n_3053_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3054 (.A1(_00490_),
    .A2(net),
    .B(n_3053_o_0),
    .C(_00884_),
    .Y(n_3054_o_0));
 OAI211xp5_ASAP7_75t_R n_3055 (.A1(n_3048_o_0),
    .A2(n_3050_o_0),
    .B(n_3051_o_0),
    .C(n_3047_o_0),
    .Y(n_3055_o_0));
 OAI21xp33_ASAP7_75t_R n_3056 (.A1(n_3047_o_0),
    .A2(n_3049_o_0),
    .B(n_3055_o_0),
    .Y(n_3056_o_0));
 NOR2xp33_ASAP7_75t_R n_3057 (.A(_00490_),
    .B(net39),
    .Y(n_3057_o_0));
 AOI211xp5_ASAP7_75t_R n_3058 (.A1(n_3056_o_0),
    .A2(net),
    .B(n_2417_o_0),
    .C(n_3057_o_0),
    .Y(n_3058_o_0));
 NOR2xp33_ASAP7_75t_R n_3059 (.A(n_3054_o_0),
    .B(n_3058_o_0),
    .Y(n_3059_o_0));
 XNOR2xp5_ASAP7_75t_R n_3060 (.A(_00996_),
    .B(_01003_),
    .Y(n_3060_o_0));
 XNOR2xp5_ASAP7_75t_R n_3061 (.A(_01116_),
    .B(n_3060_o_0),
    .Y(n_3061_o_0));
 XNOR2xp5_ASAP7_75t_R n_3062 (.A(_01036_),
    .B(_01043_),
    .Y(n_3062_o_0));
 XOR2xp5_ASAP7_75t_R n_3063 (.A(_01037_),
    .B(_01077_),
    .Y(n_3063_o_0));
 XNOR2xp5_ASAP7_75t_R n_3064 (.A(n_3062_o_0),
    .B(n_3063_o_0),
    .Y(n_3064_o_0));
 XOR2xp5_ASAP7_75t_R n_3065 (.A(_00996_),
    .B(_01003_),
    .Y(n_3065_o_0));
 NAND2xp33_ASAP7_75t_R n_3066 (.A(_01116_),
    .B(n_3065_o_0),
    .Y(n_3066_o_0));
 INVx1_ASAP7_75t_R n_3067 (.A(_01116_),
    .Y(n_3067_o_0));
 NAND2xp33_ASAP7_75t_R n_3068 (.A(n_3067_o_0),
    .B(n_3060_o_0),
    .Y(n_3068_o_0));
 NOR2xp33_ASAP7_75t_R n_3069 (.A(_01037_),
    .B(_01077_),
    .Y(n_3069_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3070 (.A1(_01037_),
    .A2(_01077_),
    .B(n_3069_o_0),
    .C(n_3062_o_0),
    .Y(n_3070_o_0));
 INVx1_ASAP7_75t_R n_3071 (.A(_01036_),
    .Y(n_3071_o_0));
 NOR2xp33_ASAP7_75t_R n_3072 (.A(_01043_),
    .B(n_3071_o_0),
    .Y(n_3072_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3073 (.A1(n_3071_o_0),
    .A2(_01043_),
    .B(n_3072_o_0),
    .C(n_3063_o_0),
    .Y(n_3073_o_0));
 AOI22xp33_ASAP7_75t_R n_3074 (.A1(n_3066_o_0),
    .A2(n_3068_o_0),
    .B1(n_3070_o_0),
    .B2(n_3073_o_0),
    .Y(n_3074_o_0));
 OAI21xp33_ASAP7_75t_R n_3075 (.A1(_00489_),
    .A2(net39),
    .B(n_2438_o_0),
    .Y(n_3075_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3076 (.A1(n_3061_o_0),
    .A2(n_3064_o_0),
    .B(n_3074_o_0),
    .C(net77),
    .D(n_3075_o_0),
    .Y(n_3076_o_0));
 NAND4xp25_ASAP7_75t_R n_3077 (.A(n_3066_o_0),
    .B(n_3068_o_0),
    .C(n_3073_o_0),
    .D(n_3070_o_0),
    .Y(n_3077_o_0));
 XOR2xp5_ASAP7_75t_R n_3078 (.A(_01036_),
    .B(_01043_),
    .Y(n_3078_o_0));
 NOR2xp33_ASAP7_75t_R n_3079 (.A(n_3078_o_0),
    .B(n_3063_o_0),
    .Y(n_3079_o_0));
 XNOR2xp5_ASAP7_75t_R n_3080 (.A(_01037_),
    .B(_01077_),
    .Y(n_3080_o_0));
 NOR2xp33_ASAP7_75t_R n_3081 (.A(n_3080_o_0),
    .B(n_3062_o_0),
    .Y(n_3081_o_0));
 NOR2xp33_ASAP7_75t_R n_3082 (.A(_01116_),
    .B(n_3065_o_0),
    .Y(n_3082_o_0));
 NOR2xp33_ASAP7_75t_R n_3083 (.A(n_3067_o_0),
    .B(n_3060_o_0),
    .Y(n_3083_o_0));
 OAI22xp33_ASAP7_75t_R n_3084 (.A1(n_3079_o_0),
    .A2(n_3081_o_0),
    .B1(n_3082_o_0),
    .B2(n_3083_o_0),
    .Y(n_3084_o_0));
 AOI211xp5_ASAP7_75t_R n_3085 (.A1(n_3077_o_0),
    .A2(n_3084_o_0),
    .B(net2),
    .C(n_2438_o_0),
    .Y(n_3085_o_0));
 NOR3xp33_ASAP7_75t_R n_3086 (.A(n_2438_o_0),
    .B(net),
    .C(_00489_),
    .Y(n_3086_o_0));
 OAI211xp5_ASAP7_75t_R n_3087 (.A1(_00490_),
    .A2(net77),
    .B(n_3053_o_0),
    .C(_00884_),
    .Y(n_3087_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3088 (.A1(n_3056_o_0),
    .A2(net77),
    .B(n_3057_o_0),
    .C(n_2417_o_0),
    .Y(n_3088_o_0));
 OAI311xp33_ASAP7_75t_R n_3089 (.A1(n_3076_o_0),
    .A2(n_3085_o_0),
    .A3(n_3086_o_0),
    .B1(n_3087_o_0),
    .C1(n_3088_o_0),
    .Y(n_3089_o_0));
 OAI21xp33_ASAP7_75t_R n_3090 (.A1(n_3060_o_0),
    .A2(n_3067_o_0),
    .B(n_3068_o_0),
    .Y(n_3090_o_0));
 OAI31xp33_ASAP7_75t_R n_3091 (.A1(n_3081_o_0),
    .A2(n_3079_o_0),
    .A3(n_3090_o_0),
    .B(n_3084_o_0),
    .Y(n_3091_o_0));
 AOI21xp33_ASAP7_75t_R n_3092 (.A1(_00489_),
    .A2(net5),
    .B(n_2438_o_0),
    .Y(n_3092_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_3093 (.A1(n_3021_o_0),
    .A2(n_3091_o_0),
    .B(n_3092_o_0),
    .C(n_3076_o_0),
    .Y(n_3093_o_0));
 OAI21xp33_ASAP7_75t_R n_3094 (.A1(n_3054_o_0),
    .A2(n_3058_o_0),
    .B(n_3093_o_0),
    .Y(n_3094_o_0));
 NAND2xp33_ASAP7_75t_R n_3095 (.A(n_3089_o_0),
    .B(n_3094_o_0),
    .Y(n_3095_o_0));
 NOR2xp33_ASAP7_75t_R n_3096 (.A(n_3045_o_0),
    .B(n_3095_o_0),
    .Y(n_3096_o_0));
 INVx1_ASAP7_75t_R n_3097 (.A(_00492_),
    .Y(n_3097_o_0));
 XOR2xp5_ASAP7_75t_R n_3098 (.A(_01038_),
    .B(n_3037_o_0),
    .Y(n_3098_o_0));
 AOI21xp33_ASAP7_75t_R n_3099 (.A1(n_3035_o_0),
    .A2(n_3098_o_0),
    .B(n_3021_o_0),
    .Y(n_3099_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3100 (.A1(n_3035_o_0),
    .A2(n_3098_o_0),
    .B(n_3099_o_0),
    .C(n_2464_o_0),
    .Y(n_3100_o_0));
 NOR2xp33_ASAP7_75t_R n_3101 (.A(n_3035_o_0),
    .B(n_3098_o_0),
    .Y(n_3101_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3102 (.A1(n_3035_o_0),
    .A2(n_3098_o_0),
    .B(n_3101_o_0),
    .C(net39),
    .D(n_3042_o_0),
    .Y(n_3102_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_3103 (.A1(n_3097_o_0),
    .A2(net39),
    .B(n_3100_o_0),
    .C(n_3102_o_0),
    .Y(n_3103_o_0));
 NOR2xp33_ASAP7_75t_R n_3104 (.A(n_3103_o_0),
    .B(n_3093_o_0),
    .Y(n_3104_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3105 (.A1(n_3032_o_0),
    .A2(net39),
    .B(n_3029_o_0),
    .C(n_2402_o_0),
    .Y(n_3105_o_0));
 OAI21x1_ASAP7_75t_R n_3106 (.A1(n_2402_o_0),
    .A2(n_3031_o_0),
    .B(n_3105_o_0),
    .Y(n_3106_o_0));
 INVx1_ASAP7_75t_R n_3107 (.A(n_3106_o_0),
    .Y(n_3107_o_0));
 NOR3xp33_ASAP7_75t_R n_3108 (.A(n_3096_o_0),
    .B(n_3104_o_0),
    .C(n_3107_o_0),
    .Y(n_3108_o_0));
 AOI31xp33_ASAP7_75t_R n_3109 (.A1(n_3034_o_0),
    .A2(net29),
    .A3(n_3059_o_0),
    .B(n_3108_o_0),
    .Y(n_3109_o_0));
 AOI21xp33_ASAP7_75t_R n_3110 (.A1(_00492_),
    .A2(net2),
    .B(n_3040_o_0),
    .Y(n_3110_o_0));
 AOI311xp33_ASAP7_75t_R n_3111 (.A1(n_3088_o_0),
    .A2(n_3087_o_0),
    .A3(n_3093_o_0),
    .B(n_3102_o_0),
    .C(n_3110_o_0),
    .Y(n_3111_o_0));
 XNOR2xp5_ASAP7_75t_R n_3112 (.A(_01039_),
    .B(_01043_),
    .Y(n_3112_o_0));
 XNOR2xp5_ASAP7_75t_R n_3113 (.A(_01080_),
    .B(_01119_),
    .Y(n_3113_o_0));
 XOR2xp5_ASAP7_75t_R n_3114 (.A(n_3112_o_0),
    .B(n_3113_o_0),
    .Y(n_3114_o_0));
 XNOR2xp5_ASAP7_75t_R n_3115 (.A(_00999_),
    .B(_01003_),
    .Y(n_3115_o_0));
 NAND2xp33_ASAP7_75t_R n_3116 (.A(_01040_),
    .B(n_3115_o_0),
    .Y(n_3116_o_0));
 OAI21xp33_ASAP7_75t_R n_3117 (.A1(_01040_),
    .A2(n_3115_o_0),
    .B(n_3116_o_0),
    .Y(n_3117_o_0));
 OAI21xp33_ASAP7_75t_R n_3118 (.A1(n_3117_o_0),
    .A2(n_3114_o_0),
    .B(net),
    .Y(n_3118_o_0));
 AOI21xp33_ASAP7_75t_R n_3119 (.A1(n_3114_o_0),
    .A2(n_3117_o_0),
    .B(n_3118_o_0),
    .Y(n_3119_o_0));
 AOI21xp33_ASAP7_75t_R n_3120 (.A1(net9),
    .A2(_00652_),
    .B(n_3119_o_0),
    .Y(n_3120_o_0));
 NAND2xp33_ASAP7_75t_R n_3121 (.A(_00888_),
    .B(n_3120_o_0),
    .Y(n_3121_o_0));
 OAI21xp33_ASAP7_75t_R n_3122 (.A1(_00888_),
    .A2(n_3120_o_0),
    .B(n_3121_o_0),
    .Y(n_3122_o_0));
 AOI21xp33_ASAP7_75t_R n_3123 (.A1(n_3111_o_0),
    .A2(n_3034_o_0),
    .B(n_3122_o_0),
    .Y(n_3123_o_0));
 INVx1_ASAP7_75t_R n_3124 (.A(n_3093_o_0),
    .Y(n_3124_o_0));
 NAND2xp5_ASAP7_75t_R n_3125 (.A(n_3088_o_0),
    .B(n_3087_o_0),
    .Y(n_3125_o_0));
 NAND2xp33_ASAP7_75t_R n_3126 (.A(n_3124_o_0),
    .B(n_3125_o_0),
    .Y(n_3126_o_0));
 NAND2xp33_ASAP7_75t_R n_3127 (.A(n_3045_o_0),
    .B(n_3126_o_0),
    .Y(n_3127_o_0));
 OAI21xp33_ASAP7_75t_R n_3128 (.A1(n_3097_o_0),
    .A2(net),
    .B(n_3100_o_0),
    .Y(n_3128_o_0));
 OA21x2_ASAP7_75t_R n_3129 (.A1(n_3058_o_0),
    .A2(n_3054_o_0),
    .B(n_3093_o_0),
    .Y(n_3129_o_0));
 AOI21xp33_ASAP7_75t_R n_3130 (.A1(n_3044_o_0),
    .A2(n_3128_o_0),
    .B(n_3129_o_0),
    .Y(n_3130_o_0));
 INVx1_ASAP7_75t_R n_3131 (.A(n_3129_o_0),
    .Y(n_3131_o_0));
 OAI21xp33_ASAP7_75t_R n_3132 (.A1(n_3045_o_0),
    .A2(n_3131_o_0),
    .B(n_3106_o_0),
    .Y(n_3132_o_0));
 XNOR2xp5_ASAP7_75t_R n_3133 (.A(_00888_),
    .B(n_3120_o_0),
    .Y(n_3133_o_0));
 OAI21xp33_ASAP7_75t_R n_3134 (.A1(n_3130_o_0),
    .A2(n_3132_o_0),
    .B(n_3133_o_0),
    .Y(n_3134_o_0));
 XOR2xp5_ASAP7_75t_R n_3135 (.A(_01001_),
    .B(_01041_),
    .Y(n_3135_o_0));
 XNOR2xp5_ASAP7_75t_R n_3136 (.A(_01042_),
    .B(_01082_),
    .Y(n_3136_o_0));
 NAND2xp33_ASAP7_75t_R n_3137 (.A(_01121_),
    .B(n_3136_o_0),
    .Y(n_3137_o_0));
 OAI21xp33_ASAP7_75t_R n_3138 (.A1(_01121_),
    .A2(n_3136_o_0),
    .B(n_3137_o_0),
    .Y(n_3138_o_0));
 NOR2xp33_ASAP7_75t_R n_3139 (.A(n_3135_o_0),
    .B(n_3138_o_0),
    .Y(n_3139_o_0));
 NOR2xp33_ASAP7_75t_R n_3140 (.A(_00650_),
    .B(net),
    .Y(n_3140_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3141 (.A1(n_3135_o_0),
    .A2(n_3138_o_0),
    .B(n_3139_o_0),
    .C(net),
    .D(n_3140_o_0),
    .Y(n_3141_o_0));
 XNOR2xp5_ASAP7_75t_R n_3142 (.A(_00890_),
    .B(n_3141_o_0),
    .Y(n_3142_o_0));
 INVx1_ASAP7_75t_R n_3143 (.A(n_3142_o_0),
    .Y(n_3143_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3144 (.A1(n_3034_o_0),
    .A2(n_3127_o_0),
    .B(n_3134_o_0),
    .C(n_3143_o_0),
    .Y(n_3144_o_0));
 NOR2xp33_ASAP7_75t_R n_3145 (.A(n_3103_o_0),
    .B(n_3034_o_0),
    .Y(n_3145_o_0));
 AOI211xp5_ASAP7_75t_R n_3146 (.A1(n_3032_o_0),
    .A2(net39),
    .B(_00887_),
    .C(n_3029_o_0),
    .Y(n_3146_o_0));
 AOI21x1_ASAP7_75t_R n_3147 (.A1(n_3031_o_0),
    .A2(_00887_),
    .B(n_3146_o_0),
    .Y(n_3147_o_0));
 AOI211xp5_ASAP7_75t_R n_3148 (.A1(n_3044_o_0),
    .A2(n_3128_o_0),
    .B(n_3059_o_0),
    .C(n_3093_o_0),
    .Y(n_3148_o_0));
 INVx1_ASAP7_75t_R n_3149 (.A(_00888_),
    .Y(n_3149_o_0));
 NAND2xp33_ASAP7_75t_R n_3150 (.A(n_3149_o_0),
    .B(n_3120_o_0),
    .Y(n_3150_o_0));
 OAI21xp33_ASAP7_75t_R n_3151 (.A1(n_3120_o_0),
    .A2(n_3149_o_0),
    .B(n_3150_o_0),
    .Y(n_3151_o_0));
 OAI31xp33_ASAP7_75t_R n_3152 (.A1(n_3147_o_0),
    .A2(n_3111_o_0),
    .A3(n_3148_o_0),
    .B(n_3151_o_0),
    .Y(n_3152_o_0));
 OAI31xp33_ASAP7_75t_R n_3153 (.A1(n_3125_o_0),
    .A2(n_3045_o_0),
    .A3(n_3124_o_0),
    .B(n_3106_o_0),
    .Y(n_3153_o_0));
 XNOR2xp5_ASAP7_75t_R n_3154 (.A(n_3149_o_0),
    .B(n_3120_o_0),
    .Y(n_3154_o_0));
 AOI31xp33_ASAP7_75t_R n_3155 (.A1(n_3045_o_0),
    .A2(n_3107_o_0),
    .A3(n_3129_o_0),
    .B(n_3154_o_0),
    .Y(n_3155_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3156 (.A1(n_3148_o_0),
    .A2(n_3153_o_0),
    .B(n_3155_o_0),
    .C(n_3143_o_0),
    .Y(n_3156_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3157 (.A1(n_3129_o_0),
    .A2(n_3145_o_0),
    .B(n_3152_o_0),
    .C(n_3156_o_0),
    .Y(n_3157_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3158 (.A1(n_3109_o_0),
    .A2(n_3123_o_0),
    .B(n_3144_o_0),
    .C(n_3157_o_0),
    .Y(n_3158_o_0));
 NOR2xp33_ASAP7_75t_R n_3159 (.A(n_3020_o_0),
    .B(n_3158_o_0),
    .Y(n_3159_o_0));
 NAND2xp33_ASAP7_75t_R n_3160 (.A(_00890_),
    .B(n_3141_o_0),
    .Y(n_3160_o_0));
 OAI21xp33_ASAP7_75t_R n_3161 (.A1(_00890_),
    .A2(n_3141_o_0),
    .B(n_3160_o_0),
    .Y(n_3161_o_0));
 AO21x1_ASAP7_75t_R n_3162 (.A1(net2),
    .A2(n_3092_o_0),
    .B(n_3085_o_0),
    .Y(n_3162_o_0));
 OAI211xp5_ASAP7_75t_R n_3163 (.A1(n_3162_o_0),
    .A2(n_3076_o_0),
    .B(n_3044_o_0),
    .C(n_3128_o_0),
    .Y(n_3163_o_0));
 NOR2xp33_ASAP7_75t_R n_3164 (.A(n_3125_o_0),
    .B(n_3163_o_0),
    .Y(n_3164_o_0));
 INVx1_ASAP7_75t_R n_3165 (.A(n_3164_o_0),
    .Y(n_3165_o_0));
 AOI22xp33_ASAP7_75t_R n_3166 (.A1(n_3094_o_0),
    .A2(n_3089_o_0),
    .B1(n_3044_o_0),
    .B2(n_3128_o_0),
    .Y(n_3166_o_0));
 NOR2xp33_ASAP7_75t_R n_3167 (.A(n_3166_o_0),
    .B(n_3107_o_0),
    .Y(n_3167_o_0));
 NOR2xp33_ASAP7_75t_R n_3168 (.A(n_3124_o_0),
    .B(n_3125_o_0),
    .Y(n_3168_o_0));
 NOR2xp33_ASAP7_75t_R n_3169 (.A(n_3103_o_0),
    .B(n_3168_o_0),
    .Y(n_3169_o_0));
 INVx1_ASAP7_75t_R n_3170 (.A(n_3169_o_0),
    .Y(n_3170_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3171 (.A1(n_3129_o_0),
    .A2(net29),
    .B(n_3170_o_0),
    .C(n_3147_o_0),
    .Y(n_3171_o_0));
 AOI21xp33_ASAP7_75t_R n_3172 (.A1(n_3165_o_0),
    .A2(n_3167_o_0),
    .B(n_3171_o_0),
    .Y(n_3172_o_0));
 NAND2xp33_ASAP7_75t_R n_3173 (.A(n_3093_o_0),
    .B(n_3125_o_0),
    .Y(n_3173_o_0));
 OAI21xp33_ASAP7_75t_R n_3174 (.A1(n_3103_o_0),
    .A2(n_3125_o_0),
    .B(n_3106_o_0),
    .Y(n_3174_o_0));
 INVx1_ASAP7_75t_R n_3175 (.A(n_3174_o_0),
    .Y(n_3175_o_0));
 NOR2xp33_ASAP7_75t_R n_3176 (.A(n_3125_o_0),
    .B(n_3045_o_0),
    .Y(n_3176_o_0));
 NOR2xp33_ASAP7_75t_R n_3177 (.A(n_3093_o_0),
    .B(n_3059_o_0),
    .Y(n_3177_o_0));
 NOR3xp33_ASAP7_75t_R n_3178 (.A(n_3176_o_0),
    .B(n_3106_o_0),
    .C(n_3177_o_0),
    .Y(n_3178_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3179 (.A1(n_3173_o_0),
    .A2(n_3175_o_0),
    .B(n_3178_o_0),
    .C(n_3133_o_0),
    .Y(n_3179_o_0));
 OAI21xp33_ASAP7_75t_R n_3180 (.A1(n_3133_o_0),
    .A2(n_3172_o_0),
    .B(n_3179_o_0),
    .Y(n_3180_o_0));
 OAI21xp33_ASAP7_75t_R n_3181 (.A1(n_3059_o_0),
    .A2(n_3163_o_0),
    .B(n_3106_o_0),
    .Y(n_3181_o_0));
 INVx1_ASAP7_75t_R n_3182 (.A(n_3181_o_0),
    .Y(n_3182_o_0));
 AOI21xp33_ASAP7_75t_R n_3183 (.A1(n_3088_o_0),
    .A2(n_3087_o_0),
    .B(n_3103_o_0),
    .Y(n_3183_o_0));
 INVx1_ASAP7_75t_R n_3184 (.A(n_3183_o_0),
    .Y(n_3184_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3185 (.A1(n_3125_o_0),
    .A2(net40),
    .B(n_3103_o_0),
    .C(n_3147_o_0),
    .Y(n_3185_o_0));
 INVx1_ASAP7_75t_R n_3186 (.A(n_3185_o_0),
    .Y(n_3186_o_0));
 OAI21xp33_ASAP7_75t_R n_3187 (.A1(n_3166_o_0),
    .A2(n_3186_o_0),
    .B(n_3133_o_0),
    .Y(n_3187_o_0));
 AOI21xp33_ASAP7_75t_R n_3188 (.A1(n_3182_o_0),
    .A2(n_3184_o_0),
    .B(n_3187_o_0),
    .Y(n_3188_o_0));
 NAND2xp33_ASAP7_75t_R n_3189 (.A(n_3125_o_0),
    .B(n_3103_o_0),
    .Y(n_3189_o_0));
 NAND2xp33_ASAP7_75t_R n_3190 (.A(n_3106_o_0),
    .B(n_3189_o_0),
    .Y(n_3190_o_0));
 NOR2xp33_ASAP7_75t_R n_3191 (.A(n_3059_o_0),
    .B(n_3163_o_0),
    .Y(n_3191_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3192 (.A1(net29),
    .A2(n_3126_o_0),
    .B(n_3147_o_0),
    .C(n_3190_o_0),
    .D(n_3191_o_0),
    .Y(n_3192_o_0));
 NOR3xp33_ASAP7_75t_R n_3193 (.A(n_3190_o_0),
    .B(n_3163_o_0),
    .C(n_3059_o_0),
    .Y(n_3193_o_0));
 OAI31xp33_ASAP7_75t_R n_3194 (.A1(n_3192_o_0),
    .A2(n_3193_o_0),
    .A3(n_3122_o_0),
    .B(n_3143_o_0),
    .Y(n_3194_o_0));
 OAI21xp33_ASAP7_75t_R n_3195 (.A1(n_3188_o_0),
    .A2(n_3194_o_0),
    .B(n_3020_o_0),
    .Y(n_3195_o_0));
 AOI21xp33_ASAP7_75t_R n_3196 (.A1(n_3161_o_0),
    .A2(n_3180_o_0),
    .B(n_3195_o_0),
    .Y(n_3196_o_0));
 NAND2xp33_ASAP7_75t_R n_3197 (.A(n_3045_o_0),
    .B(n_3106_o_0),
    .Y(n_3197_o_0));
 INVx1_ASAP7_75t_R n_3198 (.A(n_3168_o_0),
    .Y(n_3198_o_0));
 AOI211xp5_ASAP7_75t_R n_3199 (.A1(n_3103_o_0),
    .A2(n_3129_o_0),
    .B(n_3166_o_0),
    .C(n_3147_o_0),
    .Y(n_3199_o_0));
 AOI31xp33_ASAP7_75t_R n_3200 (.A1(n_3198_o_0),
    .A2(n_3106_o_0),
    .A3(net36),
    .B(n_3199_o_0),
    .Y(n_3200_o_0));
 OAI21xp33_ASAP7_75t_R n_3201 (.A1(n_3197_o_0),
    .A2(n_3129_o_0),
    .B(n_3200_o_0),
    .Y(n_3201_o_0));
 NAND2xp33_ASAP7_75t_R n_3202 (.A(n_3124_o_0),
    .B(n_3103_o_0),
    .Y(n_3202_o_0));
 OAI21xp33_ASAP7_75t_R n_3203 (.A1(n_3103_o_0),
    .A2(n_3095_o_0),
    .B(n_3106_o_0),
    .Y(n_3203_o_0));
 INVx1_ASAP7_75t_R n_3204 (.A(n_3203_o_0),
    .Y(n_3204_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3205 (.A1(n_3095_o_0),
    .A2(net36),
    .B(n_3147_o_0),
    .C(n_3133_o_0),
    .Y(n_3205_o_0));
 AOI21xp33_ASAP7_75t_R n_3206 (.A1(n_3202_o_0),
    .A2(n_3204_o_0),
    .B(n_3205_o_0),
    .Y(n_3206_o_0));
 AOI21xp33_ASAP7_75t_R n_3207 (.A1(n_3151_o_0),
    .A2(n_3201_o_0),
    .B(n_3206_o_0),
    .Y(n_3207_o_0));
 AOI21xp33_ASAP7_75t_R n_3208 (.A1(n_3125_o_0),
    .A2(n_3124_o_0),
    .B(n_3045_o_0),
    .Y(n_3208_o_0));
 NOR3xp33_ASAP7_75t_R n_3209 (.A(n_3107_o_0),
    .B(n_3208_o_0),
    .C(n_3148_o_0),
    .Y(n_3209_o_0));
 AOI211xp5_ASAP7_75t_R n_3210 (.A1(_00887_),
    .A2(n_3031_o_0),
    .B(n_3045_o_0),
    .C(n_3146_o_0),
    .Y(n_3210_o_0));
 NOR2xp33_ASAP7_75t_R n_3211 (.A(net40),
    .B(n_3103_o_0),
    .Y(n_3211_o_0));
 AOI321xp33_ASAP7_75t_R n_3212 (.A1(n_3089_o_0),
    .A2(n_3094_o_0),
    .A3(n_3210_o_0),
    .B1(n_3211_o_0),
    .B2(n_3107_o_0),
    .C(n_3154_o_0),
    .Y(n_3212_o_0));
 NAND2xp33_ASAP7_75t_R n_3213 (.A(n_3209_o_0),
    .B(n_3212_o_0),
    .Y(n_3213_o_0));
 NOR2xp33_ASAP7_75t_R n_3214 (.A(n_3125_o_0),
    .B(n_3045_o_0),
    .Y(n_3214_o_0));
 NOR2xp33_ASAP7_75t_R n_3215 (.A(n_3103_o_0),
    .B(n_3129_o_0),
    .Y(n_3215_o_0));
 OAI21xp33_ASAP7_75t_R n_3216 (.A1(n_3214_o_0),
    .A2(n_3215_o_0),
    .B(n_3107_o_0),
    .Y(n_3216_o_0));
 AOI31xp33_ASAP7_75t_R n_3217 (.A1(n_3147_o_0),
    .A2(n_3103_o_0),
    .A3(n_3129_o_0),
    .B(n_3133_o_0),
    .Y(n_3217_o_0));
 INVx1_ASAP7_75t_R n_3218 (.A(n_3208_o_0),
    .Y(n_3218_o_0));
 INVx1_ASAP7_75t_R n_3219 (.A(n_3148_o_0),
    .Y(n_3219_o_0));
 NAND3xp33_ASAP7_75t_R n_3220 (.A(n_3218_o_0),
    .B(n_3219_o_0),
    .C(n_3106_o_0),
    .Y(n_3220_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3221 (.A1(n_3216_o_0),
    .A2(n_3217_o_0),
    .B(n_3212_o_0),
    .C(n_3220_o_0),
    .Y(n_3221_o_0));
 AOI21xp33_ASAP7_75t_R n_3222 (.A1(n_3213_o_0),
    .A2(n_3221_o_0),
    .B(n_3020_o_0),
    .Y(n_3222_o_0));
 AOI21xp33_ASAP7_75t_R n_3223 (.A1(n_3020_o_0),
    .A2(n_3207_o_0),
    .B(n_3222_o_0),
    .Y(n_3223_o_0));
 NAND3xp33_ASAP7_75t_R n_3224 (.A(n_3147_o_0),
    .B(n_3045_o_0),
    .C(n_3129_o_0),
    .Y(n_3224_o_0));
 NAND2xp33_ASAP7_75t_R n_3225 (.A(n_3093_o_0),
    .B(n_3103_o_0),
    .Y(n_3225_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3226 (.A1(n_3224_o_0),
    .A2(n_3225_o_0),
    .B(n_3034_o_0),
    .C(n_3151_o_0),
    .Y(n_3226_o_0));
 NAND2xp5_ASAP7_75t_R n_3227 (.A(n_3093_o_0),
    .B(n_3045_o_0),
    .Y(n_3227_o_0));
 INVx1_ASAP7_75t_R n_3228 (.A(n_3227_o_0),
    .Y(n_3228_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3229 (.A1(n_3102_o_0),
    .A2(n_3110_o_0),
    .B(net40),
    .C(n_3125_o_0),
    .Y(n_3229_o_0));
 NAND2xp33_ASAP7_75t_R n_3230 (.A(n_3034_o_0),
    .B(n_3229_o_0),
    .Y(n_3230_o_0));
 OAI211xp5_ASAP7_75t_R n_3231 (.A1(n_3228_o_0),
    .A2(n_3181_o_0),
    .B(n_3230_o_0),
    .C(n_3133_o_0),
    .Y(n_3231_o_0));
 NOR2xp33_ASAP7_75t_R n_3232 (.A(n_3093_o_0),
    .B(n_3125_o_0),
    .Y(n_3232_o_0));
 NAND2xp33_ASAP7_75t_R n_3233 (.A(n_3034_o_0),
    .B(n_3189_o_0),
    .Y(n_3233_o_0));
 AOI211xp5_ASAP7_75t_R n_3234 (.A1(n_3232_o_0),
    .A2(net29),
    .B(n_3233_o_0),
    .C(n_3133_o_0),
    .Y(n_3234_o_0));
 AOI31xp33_ASAP7_75t_R n_3235 (.A1(n_3226_o_0),
    .A2(n_3231_o_0),
    .A3(n_3020_o_0),
    .B(n_3234_o_0),
    .Y(n_3235_o_0));
 NOR3xp33_ASAP7_75t_R n_3236 (.A(n_3126_o_0),
    .B(net29),
    .C(n_3034_o_0),
    .Y(n_3236_o_0));
 OAI211xp5_ASAP7_75t_R n_3237 (.A1(n_3102_o_0),
    .A2(n_3110_o_0),
    .B(n_3059_o_0),
    .C(n_3093_o_0),
    .Y(n_3237_o_0));
 INVx1_ASAP7_75t_R n_3238 (.A(n_3146_o_0),
    .Y(n_3238_o_0));
 AO21x1_ASAP7_75t_R n_3239 (.A1(n_3238_o_0),
    .A2(n_3033_o_0),
    .B(n_3166_o_0),
    .Y(n_3239_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3240 (.A1(n_3034_o_0),
    .A2(n_3237_o_0),
    .B(n_3239_o_0),
    .C(n_3151_o_0),
    .Y(n_3240_o_0));
 INVx1_ASAP7_75t_R n_3241 (.A(n_3020_o_0),
    .Y(n_3241_o_0));
 OAI21xp33_ASAP7_75t_R n_3242 (.A1(n_3236_o_0),
    .A2(n_3240_o_0),
    .B(n_3241_o_0),
    .Y(n_3242_o_0));
 NAND3xp33_ASAP7_75t_R n_3243 (.A(n_3235_o_0),
    .B(n_3242_o_0),
    .C(n_3143_o_0),
    .Y(n_3243_o_0));
 NAND2xp33_ASAP7_75t_R n_3244 (.A(_00889_),
    .B(n_3009_o_0),
    .Y(n_3244_o_0));
 OAI21xp5_ASAP7_75t_R n_3245 (.A1(_00889_),
    .A2(n_3009_o_0),
    .B(n_3244_o_0),
    .Y(n_3245_o_0));
 OAI211xp5_ASAP7_75t_R n_3246 (.A1(n_3223_o_0),
    .A2(n_3143_o_0),
    .B(n_3243_o_0),
    .C(n_3245_o_0),
    .Y(n_3246_o_0));
 OAI31xp33_ASAP7_75t_R n_3247 (.A1(n_3010_o_0),
    .A2(n_3159_o_0),
    .A3(n_3196_o_0),
    .B(n_3246_o_0),
    .Y(n_3247_o_0));
 OAI21xp33_ASAP7_75t_R n_3248 (.A1(n_3059_o_0),
    .A2(n_3093_o_0),
    .B(n_3045_o_0),
    .Y(n_3248_o_0));
 AOI21xp33_ASAP7_75t_R n_3249 (.A1(n_3093_o_0),
    .A2(n_3103_o_0),
    .B(n_3106_o_0),
    .Y(n_3249_o_0));
 NAND2xp33_ASAP7_75t_R n_3250 (.A(n_3248_o_0),
    .B(n_3249_o_0),
    .Y(n_3250_o_0));
 NAND2xp33_ASAP7_75t_R n_3251 (.A(n_3202_o_0),
    .B(n_3175_o_0),
    .Y(n_3251_o_0));
 INVx1_ASAP7_75t_R n_3252 (.A(n_3132_o_0),
    .Y(n_3252_o_0));
 NOR2xp33_ASAP7_75t_R n_3253 (.A(n_3093_o_0),
    .B(n_3059_o_0),
    .Y(n_3253_o_0));
 NOR3xp33_ASAP7_75t_R n_3254 (.A(n_3253_o_0),
    .B(n_3045_o_0),
    .C(n_3147_o_0),
    .Y(n_3254_o_0));
 AOI21xp33_ASAP7_75t_R n_3255 (.A1(n_3184_o_0),
    .A2(n_3227_o_0),
    .B(n_3106_o_0),
    .Y(n_3255_o_0));
 AOI211xp5_ASAP7_75t_R n_3256 (.A1(n_3252_o_0),
    .A2(n_3184_o_0),
    .B(n_3254_o_0),
    .C(n_3255_o_0),
    .Y(n_3256_o_0));
 INVx1_ASAP7_75t_R n_3257 (.A(n_3010_o_0),
    .Y(n_3257_o_0));
 AOI32xp33_ASAP7_75t_R n_3258 (.A1(n_3245_o_0),
    .A2(n_3250_o_0),
    .A3(n_3251_o_0),
    .B1(n_3256_o_0),
    .B2(n_3257_o_0),
    .Y(n_3258_o_0));
 INVx1_ASAP7_75t_R n_3259 (.A(n_3232_o_0),
    .Y(n_3259_o_0));
 INVx1_ASAP7_75t_R n_3260 (.A(n_3153_o_0),
    .Y(n_3260_o_0));
 OAI21xp33_ASAP7_75t_R n_3261 (.A1(net36),
    .A2(n_3259_o_0),
    .B(n_3260_o_0),
    .Y(n_3261_o_0));
 NAND2xp33_ASAP7_75t_R n_3262 (.A(net40),
    .B(net36),
    .Y(n_3262_o_0));
 NAND3xp33_ASAP7_75t_R n_3263 (.A(n_3245_o_0),
    .B(n_3262_o_0),
    .C(n_3034_o_0),
    .Y(n_3263_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3264 (.A1(n_3261_o_0),
    .A2(n_3263_o_0),
    .B(n_3133_o_0),
    .C(n_3142_o_0),
    .Y(n_3264_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3265 (.A1(n_3258_o_0),
    .A2(n_3133_o_0),
    .B(n_3264_o_0),
    .C(n_3020_o_0),
    .Y(n_3265_o_0));
 AOI21xp33_ASAP7_75t_R n_3266 (.A1(n_3045_o_0),
    .A2(n_3232_o_0),
    .B(n_3107_o_0),
    .Y(n_3266_o_0));
 NAND2xp33_ASAP7_75t_R n_3267 (.A(n_3189_o_0),
    .B(n_3266_o_0),
    .Y(n_3267_o_0));
 NOR2xp33_ASAP7_75t_R n_3268 (.A(n_3045_o_0),
    .B(n_3131_o_0),
    .Y(n_3268_o_0));
 INVx1_ASAP7_75t_R n_3269 (.A(n_3245_o_0),
    .Y(n_3269_o_0));
 OA211x2_ASAP7_75t_R n_3270 (.A1(n_3268_o_0),
    .A2(n_3174_o_0),
    .B(n_3250_o_0),
    .C(n_3269_o_0),
    .Y(n_3270_o_0));
 AOI31xp33_ASAP7_75t_R n_3271 (.A1(n_3239_o_0),
    .A2(n_3245_o_0),
    .A3(n_3267_o_0),
    .B(n_3270_o_0),
    .Y(n_3271_o_0));
 AOI31xp33_ASAP7_75t_R n_3272 (.A1(n_3089_o_0),
    .A2(n_3045_o_0),
    .A3(n_3094_o_0),
    .B(n_3147_o_0),
    .Y(n_3272_o_0));
 OAI21xp33_ASAP7_75t_R n_3273 (.A1(n_3129_o_0),
    .A2(n_3045_o_0),
    .B(n_3106_o_0),
    .Y(n_3273_o_0));
 NOR2xp33_ASAP7_75t_R n_3274 (.A(n_3093_o_0),
    .B(n_3125_o_0),
    .Y(n_3274_o_0));
 AOI21xp33_ASAP7_75t_R n_3275 (.A1(n_3044_o_0),
    .A2(n_3128_o_0),
    .B(n_3274_o_0),
    .Y(n_3275_o_0));
 NOR2xp33_ASAP7_75t_R n_3276 (.A(n_3273_o_0),
    .B(n_3275_o_0),
    .Y(n_3276_o_0));
 AOI21xp33_ASAP7_75t_R n_3277 (.A1(n_3165_o_0),
    .A2(n_3272_o_0),
    .B(n_3276_o_0),
    .Y(n_3277_o_0));
 INVx1_ASAP7_75t_R n_3278 (.A(n_3214_o_0),
    .Y(n_3278_o_0));
 OAI21xp33_ASAP7_75t_R n_3279 (.A1(n_3034_o_0),
    .A2(n_3278_o_0),
    .B(n_3257_o_0),
    .Y(n_3279_o_0));
 INVx1_ASAP7_75t_R n_3280 (.A(n_3215_o_0),
    .Y(n_3280_o_0));
 INVx1_ASAP7_75t_R n_3281 (.A(n_3095_o_0),
    .Y(n_3281_o_0));
 NAND3xp33_ASAP7_75t_R n_3282 (.A(n_3281_o_0),
    .B(n_3107_o_0),
    .C(n_3103_o_0),
    .Y(n_3282_o_0));
 OAI211xp5_ASAP7_75t_R n_3283 (.A1(n_3106_o_0),
    .A2(n_3280_o_0),
    .B(n_3282_o_0),
    .C(n_3224_o_0),
    .Y(n_3283_o_0));
 OAI21xp33_ASAP7_75t_R n_3284 (.A1(n_3279_o_0),
    .A2(n_3283_o_0),
    .B(n_3133_o_0),
    .Y(n_3284_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3285 (.A1(n_3245_o_0),
    .A2(n_3277_o_0),
    .B(n_3284_o_0),
    .C(n_3143_o_0),
    .Y(n_3285_o_0));
 AOI21xp33_ASAP7_75t_R n_3286 (.A1(n_3154_o_0),
    .A2(n_3271_o_0),
    .B(n_3285_o_0),
    .Y(n_3286_o_0));
 INVx1_ASAP7_75t_R n_3287 (.A(n_3104_o_0),
    .Y(n_3287_o_0));
 NOR3xp33_ASAP7_75t_R n_3288 (.A(n_3253_o_0),
    .B(net29),
    .C(n_3147_o_0),
    .Y(n_3288_o_0));
 AOI31xp33_ASAP7_75t_R n_3289 (.A1(n_3106_o_0),
    .A2(n_3287_o_0),
    .A3(n_3173_o_0),
    .B(n_3288_o_0),
    .Y(n_3289_o_0));
 NOR2xp33_ASAP7_75t_R n_3290 (.A(n_3147_o_0),
    .B(n_3166_o_0),
    .Y(n_3290_o_0));
 AOI21xp33_ASAP7_75t_R n_3291 (.A1(n_3045_o_0),
    .A2(n_3126_o_0),
    .B(n_3107_o_0),
    .Y(n_3291_o_0));
 AO21x1_ASAP7_75t_R n_3292 (.A1(n_3291_o_0),
    .A2(n_3278_o_0),
    .B(n_3151_o_0),
    .Y(n_3292_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3293 (.A1(n_3189_o_0),
    .A2(n_3290_o_0),
    .B(n_3292_o_0),
    .C(n_3257_o_0),
    .Y(n_3293_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3294 (.A1(n_3154_o_0),
    .A2(n_3289_o_0),
    .B(n_3293_o_0),
    .C(n_3142_o_0),
    .Y(n_3294_o_0));
 AOI211xp5_ASAP7_75t_R n_3295 (.A1(n_3107_o_0),
    .A2(n_3163_o_0),
    .B(n_3236_o_0),
    .C(n_3154_o_0),
    .Y(n_3295_o_0));
 NAND2xp33_ASAP7_75t_R n_3296 (.A(n_3103_o_0),
    .B(n_3095_o_0),
    .Y(n_3296_o_0));
 INVx1_ASAP7_75t_R n_3297 (.A(n_3296_o_0),
    .Y(n_3297_o_0));
 OAI31xp33_ASAP7_75t_R n_3298 (.A1(n_3147_o_0),
    .A2(n_3297_o_0),
    .A3(n_3275_o_0),
    .B(n_3154_o_0),
    .Y(n_3298_o_0));
 OAI21xp33_ASAP7_75t_R n_3299 (.A1(n_3209_o_0),
    .A2(n_3298_o_0),
    .B(n_3010_o_0),
    .Y(n_3299_o_0));
 AOI21xp33_ASAP7_75t_R n_3300 (.A1(n_3227_o_0),
    .A2(n_3295_o_0),
    .B(n_3299_o_0),
    .Y(n_3300_o_0));
 INVx1_ASAP7_75t_R n_3301 (.A(n_3126_o_0),
    .Y(n_3301_o_0));
 AOI211xp5_ASAP7_75t_R n_3302 (.A1(n_3301_o_0),
    .A2(net36),
    .B(n_3147_o_0),
    .C(n_3166_o_0),
    .Y(n_3302_o_0));
 AOI31xp33_ASAP7_75t_R n_3303 (.A1(n_3106_o_0),
    .A2(n_3278_o_0),
    .A3(n_3280_o_0),
    .B(n_3302_o_0),
    .Y(n_3303_o_0));
 AOI21xp33_ASAP7_75t_R n_3304 (.A1(n_3227_o_0),
    .A2(n_3185_o_0),
    .B(n_3245_o_0),
    .Y(n_3304_o_0));
 OAI21xp33_ASAP7_75t_R n_3305 (.A1(n_3197_o_0),
    .A2(n_3232_o_0),
    .B(n_3304_o_0),
    .Y(n_3305_o_0));
 OAI21xp33_ASAP7_75t_R n_3306 (.A1(n_3269_o_0),
    .A2(n_3303_o_0),
    .B(n_3305_o_0),
    .Y(n_3306_o_0));
 OAI21xp33_ASAP7_75t_R n_3307 (.A1(n_3183_o_0),
    .A2(n_3232_o_0),
    .B(n_3107_o_0),
    .Y(n_3307_o_0));
 AOI31xp33_ASAP7_75t_R n_3308 (.A1(n_3089_o_0),
    .A2(n_3103_o_0),
    .A3(n_3094_o_0),
    .B(n_3034_o_0),
    .Y(n_3308_o_0));
 OAI21xp33_ASAP7_75t_R n_3309 (.A1(n_3059_o_0),
    .A2(net36),
    .B(n_3308_o_0),
    .Y(n_3309_o_0));
 NAND3xp33_ASAP7_75t_R n_3310 (.A(n_3307_o_0),
    .B(n_3309_o_0),
    .C(n_3245_o_0),
    .Y(n_3310_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3311 (.A1(n_3163_o_0),
    .A2(n_3125_o_0),
    .B(n_3272_o_0),
    .C(n_3010_o_0),
    .Y(n_3311_o_0));
 OAI31xp33_ASAP7_75t_R n_3312 (.A1(n_3034_o_0),
    .A2(n_3126_o_0),
    .A3(net36),
    .B(n_3311_o_0),
    .Y(n_3312_o_0));
 AOI31xp33_ASAP7_75t_R n_3313 (.A1(n_3154_o_0),
    .A2(n_3310_o_0),
    .A3(n_3312_o_0),
    .B(n_3142_o_0),
    .Y(n_3313_o_0));
 OAI21xp33_ASAP7_75t_R n_3314 (.A1(n_3151_o_0),
    .A2(n_3306_o_0),
    .B(n_3313_o_0),
    .Y(n_3314_o_0));
 OAI21xp33_ASAP7_75t_R n_3315 (.A1(n_3294_o_0),
    .A2(n_3300_o_0),
    .B(n_3314_o_0),
    .Y(n_3315_o_0));
 OAI22xp33_ASAP7_75t_R n_3316 (.A1(n_3265_o_0),
    .A2(n_3286_o_0),
    .B1(n_3315_o_0),
    .B2(n_3020_o_0),
    .Y(n_3316_o_0));
 OAI211xp5_ASAP7_75t_R n_3317 (.A1(n_3125_o_0),
    .A2(n_3045_o_0),
    .B(n_3106_o_0),
    .C(net40),
    .Y(n_3317_o_0));
 OAI31xp33_ASAP7_75t_R n_3318 (.A1(n_3147_o_0),
    .A2(n_3169_o_0),
    .A3(n_3096_o_0),
    .B(n_3317_o_0),
    .Y(n_3318_o_0));
 NAND2xp33_ASAP7_75t_R n_3319 (.A(n_3034_o_0),
    .B(n_3173_o_0),
    .Y(n_3319_o_0));
 OAI21xp33_ASAP7_75t_R n_3320 (.A1(n_3319_o_0),
    .A2(n_3104_o_0),
    .B(n_3154_o_0),
    .Y(n_3320_o_0));
 AOI21xp33_ASAP7_75t_R n_3321 (.A1(n_3106_o_0),
    .A2(n_3262_o_0),
    .B(n_3320_o_0),
    .Y(n_3321_o_0));
 AOI21xp33_ASAP7_75t_R n_3322 (.A1(n_3122_o_0),
    .A2(n_3318_o_0),
    .B(n_3321_o_0),
    .Y(n_3322_o_0));
 AOI31xp33_ASAP7_75t_R n_3323 (.A1(n_3034_o_0),
    .A2(n_3296_o_0),
    .A3(n_3219_o_0),
    .B(n_3122_o_0),
    .Y(n_3323_o_0));
 OAI31xp33_ASAP7_75t_R n_3324 (.A1(net40),
    .A2(net36),
    .A3(n_3107_o_0),
    .B(n_3323_o_0),
    .Y(n_3324_o_0));
 AOI31xp33_ASAP7_75t_R n_3325 (.A1(n_3034_o_0),
    .A2(n_3184_o_0),
    .A3(n_3225_o_0),
    .B(n_3151_o_0),
    .Y(n_3325_o_0));
 OAI31xp33_ASAP7_75t_R n_3326 (.A1(n_3096_o_0),
    .A2(n_3107_o_0),
    .A3(n_3104_o_0),
    .B(n_3325_o_0),
    .Y(n_3326_o_0));
 AND3x1_ASAP7_75t_R n_3327 (.A(n_3324_o_0),
    .B(n_3326_o_0),
    .C(n_3257_o_0),
    .Y(n_3327_o_0));
 AOI211xp5_ASAP7_75t_R n_3328 (.A1(n_3322_o_0),
    .A2(n_3245_o_0),
    .B(n_3327_o_0),
    .C(n_3161_o_0),
    .Y(n_3328_o_0));
 OAI21xp33_ASAP7_75t_R n_3329 (.A1(n_3103_o_0),
    .A2(n_3125_o_0),
    .B(n_3034_o_0),
    .Y(n_3329_o_0));
 OA21x2_ASAP7_75t_R n_3330 (.A1(n_3164_o_0),
    .A2(n_3329_o_0),
    .B(n_3133_o_0),
    .Y(n_3330_o_0));
 INVx1_ASAP7_75t_R n_3331 (.A(n_3197_o_0),
    .Y(n_3331_o_0));
 OAI21xp33_ASAP7_75t_R n_3332 (.A1(n_3208_o_0),
    .A2(n_3239_o_0),
    .B(n_3154_o_0),
    .Y(n_3332_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3333 (.A1(n_3131_o_0),
    .A2(n_3331_o_0),
    .B(n_3332_o_0),
    .C(n_3257_o_0),
    .Y(n_3333_o_0));
 OAI21xp33_ASAP7_75t_R n_3334 (.A1(n_3147_o_0),
    .A2(n_3211_o_0),
    .B(n_3181_o_0),
    .Y(n_3334_o_0));
 NAND3xp33_ASAP7_75t_R n_3335 (.A(n_3147_o_0),
    .B(n_3124_o_0),
    .C(net36),
    .Y(n_3335_o_0));
 OAI211xp5_ASAP7_75t_R n_3336 (.A1(n_3059_o_0),
    .A2(n_3163_o_0),
    .B(n_3287_o_0),
    .C(n_3034_o_0),
    .Y(n_3336_o_0));
 AOI31xp33_ASAP7_75t_R n_3337 (.A1(n_3335_o_0),
    .A2(n_3336_o_0),
    .A3(n_3133_o_0),
    .B(n_3269_o_0),
    .Y(n_3337_o_0));
 OAI21xp33_ASAP7_75t_R n_3338 (.A1(n_3122_o_0),
    .A2(n_3334_o_0),
    .B(n_3337_o_0),
    .Y(n_3338_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3339 (.A1(n_3261_o_0),
    .A2(n_3330_o_0),
    .B(n_3333_o_0),
    .C(n_3338_o_0),
    .Y(n_3339_o_0));
 NOR2xp33_ASAP7_75t_R n_3340 (.A(n_3143_o_0),
    .B(n_3339_o_0),
    .Y(n_3340_o_0));
 INVx1_ASAP7_75t_R n_3341 (.A(n_3291_o_0),
    .Y(n_3341_o_0));
 AOI21xp33_ASAP7_75t_R n_3342 (.A1(n_3059_o_0),
    .A2(n_3124_o_0),
    .B(n_3045_o_0),
    .Y(n_3342_o_0));
 OA21x2_ASAP7_75t_R n_3343 (.A1(n_3341_o_0),
    .A2(n_3342_o_0),
    .B(n_3336_o_0),
    .Y(n_3343_o_0));
 OAI31xp33_ASAP7_75t_R n_3344 (.A1(n_3154_o_0),
    .A2(n_3343_o_0),
    .A3(n_3269_o_0),
    .B(n_3142_o_0),
    .Y(n_3344_o_0));
 AOI21xp33_ASAP7_75t_R n_3345 (.A1(n_3219_o_0),
    .A2(n_3218_o_0),
    .B(n_3106_o_0),
    .Y(n_3345_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3346 (.A1(net40),
    .A2(net36),
    .B(n_3308_o_0),
    .C(n_3345_o_0),
    .Y(n_3346_o_0));
 AND3x1_ASAP7_75t_R n_3347 (.A(n_3346_o_0),
    .B(n_3245_o_0),
    .C(n_3151_o_0),
    .Y(n_3347_o_0));
 NOR2xp33_ASAP7_75t_R n_3348 (.A(n_3125_o_0),
    .B(n_3103_o_0),
    .Y(n_3348_o_0));
 OAI211xp5_ASAP7_75t_R n_3349 (.A1(n_3095_o_0),
    .A2(net36),
    .B(n_3225_o_0),
    .C(n_3106_o_0),
    .Y(n_3349_o_0));
 OAI31xp33_ASAP7_75t_R n_3350 (.A1(n_3147_o_0),
    .A2(n_3268_o_0),
    .A3(n_3348_o_0),
    .B(n_3349_o_0),
    .Y(n_3350_o_0));
 OAI31xp33_ASAP7_75t_R n_3351 (.A1(n_3275_o_0),
    .A2(n_3164_o_0),
    .A3(n_3147_o_0),
    .B(n_3181_o_0),
    .Y(n_3351_o_0));
 OAI21xp33_ASAP7_75t_R n_3352 (.A1(n_3122_o_0),
    .A2(n_3351_o_0),
    .B(n_3257_o_0),
    .Y(n_3352_o_0));
 AOI21xp33_ASAP7_75t_R n_3353 (.A1(n_3133_o_0),
    .A2(n_3350_o_0),
    .B(n_3352_o_0),
    .Y(n_3353_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3354 (.A1(n_3168_o_0),
    .A2(net36),
    .B(n_3174_o_0),
    .C(n_3154_o_0),
    .Y(n_3354_o_0));
 AO21x1_ASAP7_75t_R n_3355 (.A1(n_3296_o_0),
    .A2(n_3272_o_0),
    .B(n_3354_o_0),
    .Y(n_3355_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3356 (.A1(n_3102_o_0),
    .A2(n_3110_o_0),
    .B(n_3168_o_0),
    .C(n_3147_o_0),
    .Y(n_3356_o_0));
 OAI31xp33_ASAP7_75t_R n_3357 (.A1(n_3045_o_0),
    .A2(net40),
    .A3(n_3125_o_0),
    .B(n_3106_o_0),
    .Y(n_3357_o_0));
 OAI21xp33_ASAP7_75t_R n_3358 (.A1(n_3348_o_0),
    .A2(n_3357_o_0),
    .B(n_3133_o_0),
    .Y(n_3358_o_0));
 AO21x1_ASAP7_75t_R n_3359 (.A1(n_3356_o_0),
    .A2(n_3225_o_0),
    .B(n_3358_o_0),
    .Y(n_3359_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3360 (.A1(n_3034_o_0),
    .A2(n_3124_o_0),
    .B(net36),
    .C(n_3151_o_0),
    .Y(n_3360_o_0));
 INVx1_ASAP7_75t_R n_3361 (.A(n_3237_o_0),
    .Y(n_3361_o_0));
 AOI22xp33_ASAP7_75t_R n_3362 (.A1(n_3361_o_0),
    .A2(n_3147_o_0),
    .B1(n_3133_o_0),
    .B2(n_3357_o_0),
    .Y(n_3362_o_0));
 AOI211xp5_ASAP7_75t_R n_3363 (.A1(n_3301_o_0),
    .A2(n_3103_o_0),
    .B(n_3147_o_0),
    .C(n_3348_o_0),
    .Y(n_3363_o_0));
 OA221x2_ASAP7_75t_R n_3364 (.A1(n_3208_o_0),
    .A2(n_3360_o_0),
    .B1(n_3362_o_0),
    .B2(n_3363_o_0),
    .C(n_3245_o_0),
    .Y(n_3364_o_0));
 AOI31xp33_ASAP7_75t_R n_3365 (.A1(n_3257_o_0),
    .A2(n_3355_o_0),
    .A3(n_3359_o_0),
    .B(n_3364_o_0),
    .Y(n_3365_o_0));
 OAI321xp33_ASAP7_75t_R n_3366 (.A1(n_3344_o_0),
    .A2(n_3347_o_0),
    .A3(n_3353_o_0),
    .B1(n_3142_o_0),
    .B2(n_3365_o_0),
    .C(n_3020_o_0),
    .Y(n_3366_o_0));
 OAI31xp33_ASAP7_75t_R n_3367 (.A1(n_3020_o_0),
    .A2(n_3328_o_0),
    .A3(n_3340_o_0),
    .B(n_3366_o_0),
    .Y(n_3367_o_0));
 OAI31xp33_ASAP7_75t_R n_3368 (.A1(n_3147_o_0),
    .A2(n_3275_o_0),
    .A3(n_3208_o_0),
    .B(n_3349_o_0),
    .Y(n_3368_o_0));
 NOR2xp33_ASAP7_75t_R n_3369 (.A(n_3122_o_0),
    .B(n_3368_o_0),
    .Y(n_3369_o_0));
 AOI211xp5_ASAP7_75t_R n_3370 (.A1(n_3095_o_0),
    .A2(n_3103_o_0),
    .B(n_3215_o_0),
    .C(n_3147_o_0),
    .Y(n_3370_o_0));
 AOI31xp33_ASAP7_75t_R n_3371 (.A1(n_3106_o_0),
    .A2(n_3170_o_0),
    .A3(n_3278_o_0),
    .B(n_3370_o_0),
    .Y(n_3371_o_0));
 OAI21xp33_ASAP7_75t_R n_3372 (.A1(n_3154_o_0),
    .A2(n_3371_o_0),
    .B(n_3269_o_0),
    .Y(n_3372_o_0));
 INVx1_ASAP7_75t_R n_3373 (.A(n_3225_o_0),
    .Y(n_3373_o_0));
 NOR3xp33_ASAP7_75t_R n_3374 (.A(n_3373_o_0),
    .B(n_3183_o_0),
    .C(n_3107_o_0),
    .Y(n_3374_o_0));
 AOI21xp33_ASAP7_75t_R n_3375 (.A1(n_3225_o_0),
    .A2(n_3290_o_0),
    .B(n_3122_o_0),
    .Y(n_3375_o_0));
 OAI21xp33_ASAP7_75t_R n_3376 (.A1(n_3174_o_0),
    .A2(n_3253_o_0),
    .B(n_3375_o_0),
    .Y(n_3376_o_0));
 OAI211xp5_ASAP7_75t_R n_3377 (.A1(n_3205_o_0),
    .A2(n_3374_o_0),
    .B(n_3376_o_0),
    .C(n_3245_o_0),
    .Y(n_3377_o_0));
 OAI21xp33_ASAP7_75t_R n_3378 (.A1(n_3369_o_0),
    .A2(n_3372_o_0),
    .B(n_3377_o_0),
    .Y(n_3378_o_0));
 OA21x2_ASAP7_75t_R n_3379 (.A1(net36),
    .A2(n_3232_o_0),
    .B(n_3308_o_0),
    .Y(n_3379_o_0));
 INVx1_ASAP7_75t_R n_3380 (.A(n_3249_o_0),
    .Y(n_3380_o_0));
 OAI31xp33_ASAP7_75t_R n_3381 (.A1(n_3169_o_0),
    .A2(n_3380_o_0),
    .A3(n_3176_o_0),
    .B(n_3151_o_0),
    .Y(n_3381_o_0));
 INVx1_ASAP7_75t_R n_3382 (.A(n_3111_o_0),
    .Y(n_3382_o_0));
 AOI21xp33_ASAP7_75t_R n_3383 (.A1(n_3382_o_0),
    .A2(n_3167_o_0),
    .B(n_3178_o_0),
    .Y(n_3383_o_0));
 AOI21xp33_ASAP7_75t_R n_3384 (.A1(n_3122_o_0),
    .A2(n_3383_o_0),
    .B(n_3245_o_0),
    .Y(n_3384_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3385 (.A1(n_3059_o_0),
    .A2(n_3163_o_0),
    .B(n_3034_o_0),
    .C(n_3122_o_0),
    .Y(n_3385_o_0));
 OAI21xp33_ASAP7_75t_R n_3386 (.A1(n_3174_o_0),
    .A2(n_3253_o_0),
    .B(n_3385_o_0),
    .Y(n_3386_o_0));
 AOI21xp33_ASAP7_75t_R n_3387 (.A1(n_3059_o_0),
    .A2(n_3093_o_0),
    .B(n_3045_o_0),
    .Y(n_3387_o_0));
 AOI21xp33_ASAP7_75t_R n_3388 (.A1(n_3227_o_0),
    .A2(n_3185_o_0),
    .B(n_3151_o_0),
    .Y(n_3388_o_0));
 OAI21xp33_ASAP7_75t_R n_3389 (.A1(n_3203_o_0),
    .A2(n_3387_o_0),
    .B(n_3388_o_0),
    .Y(n_3389_o_0));
 AOI21xp33_ASAP7_75t_R n_3390 (.A1(n_3386_o_0),
    .A2(n_3389_o_0),
    .B(n_3257_o_0),
    .Y(n_3390_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3391 (.A1(n_3379_o_0),
    .A2(n_3381_o_0),
    .B(n_3384_o_0),
    .C(n_3390_o_0),
    .Y(n_3391_o_0));
 AOI22xp33_ASAP7_75t_R n_3392 (.A1(n_3378_o_0),
    .A2(n_3161_o_0),
    .B1(n_3143_o_0),
    .B2(n_3391_o_0),
    .Y(n_3392_o_0));
 NAND3xp33_ASAP7_75t_R n_3393 (.A(n_3287_o_0),
    .B(n_3173_o_0),
    .C(n_3106_o_0),
    .Y(n_3393_o_0));
 INVx1_ASAP7_75t_R n_3394 (.A(n_3342_o_0),
    .Y(n_3394_o_0));
 AOI21xp33_ASAP7_75t_R n_3395 (.A1(n_3237_o_0),
    .A2(n_3189_o_0),
    .B(n_3106_o_0),
    .Y(n_3395_o_0));
 AOI211xp5_ASAP7_75t_R n_3396 (.A1(n_3167_o_0),
    .A2(n_3394_o_0),
    .B(n_3151_o_0),
    .C(n_3395_o_0),
    .Y(n_3396_o_0));
 AOI31xp33_ASAP7_75t_R n_3397 (.A1(n_3151_o_0),
    .A2(n_3216_o_0),
    .A3(n_3393_o_0),
    .B(n_3396_o_0),
    .Y(n_3397_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3398 (.A1(net29),
    .A2(n_3232_o_0),
    .B(n_3153_o_0),
    .C(n_3329_o_0),
    .D(n_3387_o_0),
    .Y(n_3398_o_0));
 NOR3xp33_ASAP7_75t_R n_3399 (.A(n_3153_o_0),
    .B(net29),
    .C(n_3168_o_0),
    .Y(n_3399_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3400 (.A1(n_3398_o_0),
    .A2(n_3399_o_0),
    .B(n_3151_o_0),
    .C(n_3257_o_0),
    .Y(n_3400_o_0));
 AOI21xp33_ASAP7_75t_R n_3401 (.A1(n_3358_o_0),
    .A2(n_3400_o_0),
    .B(n_3161_o_0),
    .Y(n_3401_o_0));
 OAI21xp33_ASAP7_75t_R n_3402 (.A1(n_3010_o_0),
    .A2(n_3397_o_0),
    .B(n_3401_o_0),
    .Y(n_3402_o_0));
 NOR2xp33_ASAP7_75t_R n_3403 (.A(net29),
    .B(n_3147_o_0),
    .Y(n_3403_o_0));
 OAI21xp33_ASAP7_75t_R n_3404 (.A1(n_3104_o_0),
    .A2(n_3153_o_0),
    .B(n_3155_o_0),
    .Y(n_3404_o_0));
 OAI21xp33_ASAP7_75t_R n_3405 (.A1(n_3342_o_0),
    .A2(n_3329_o_0),
    .B(n_3154_o_0),
    .Y(n_3405_o_0));
 AOI211xp5_ASAP7_75t_R n_3406 (.A1(n_3167_o_0),
    .A2(n_3189_o_0),
    .B(n_3405_o_0),
    .C(n_3257_o_0),
    .Y(n_3406_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3407 (.A1(n_3403_o_0),
    .A2(n_3095_o_0),
    .B(n_3404_o_0),
    .C(n_3406_o_0),
    .Y(n_3407_o_0));
 NOR3xp33_ASAP7_75t_R n_3408 (.A(n_3131_o_0),
    .B(n_3106_o_0),
    .C(n_3103_o_0),
    .Y(n_3408_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3409 (.A1(n_3147_o_0),
    .A2(n_3166_o_0),
    .B(n_3408_o_0),
    .C(n_3133_o_0),
    .Y(n_3409_o_0));
 OAI211xp5_ASAP7_75t_R n_3410 (.A1(n_3354_o_0),
    .A2(n_3356_o_0),
    .B(n_3409_o_0),
    .C(n_3257_o_0),
    .Y(n_3410_o_0));
 AOI211xp5_ASAP7_75t_R n_3411 (.A1(n_3260_o_0),
    .A2(n_3287_o_0),
    .B(n_3154_o_0),
    .C(n_3408_o_0),
    .Y(n_3411_o_0));
 OAI311xp33_ASAP7_75t_R n_3412 (.A1(net29),
    .A2(n_3281_o_0),
    .A3(n_3147_o_0),
    .B1(n_3010_o_0),
    .C1(n_3411_o_0),
    .Y(n_3412_o_0));
 NAND4xp25_ASAP7_75t_R n_3413 (.A(n_3407_o_0),
    .B(n_3410_o_0),
    .C(n_3412_o_0),
    .D(n_3142_o_0),
    .Y(n_3413_o_0));
 AO21x1_ASAP7_75t_R n_3414 (.A1(n_3402_o_0),
    .A2(n_3413_o_0),
    .B(n_3241_o_0),
    .Y(n_3414_o_0));
 OAI21xp33_ASAP7_75t_R n_3415 (.A1(n_3020_o_0),
    .A2(n_3392_o_0),
    .B(n_3414_o_0),
    .Y(n_3415_o_0));
 AOI21xp33_ASAP7_75t_R n_3416 (.A1(n_3202_o_0),
    .A2(n_3280_o_0),
    .B(n_3106_o_0),
    .Y(n_3416_o_0));
 NOR3xp33_ASAP7_75t_R n_3417 (.A(n_3416_o_0),
    .B(n_3209_o_0),
    .C(n_3133_o_0),
    .Y(n_3417_o_0));
 OAI32xp33_ASAP7_75t_R n_3418 (.A1(n_3147_o_0),
    .A2(n_3148_o_0),
    .A3(n_3373_o_0),
    .B1(n_3341_o_0),
    .B2(n_3342_o_0),
    .Y(n_3418_o_0));
 OAI21xp33_ASAP7_75t_R n_3419 (.A1(n_3154_o_0),
    .A2(n_3418_o_0),
    .B(n_3010_o_0),
    .Y(n_3419_o_0));
 NOR3xp33_ASAP7_75t_R n_3420 (.A(n_3297_o_0),
    .B(n_3275_o_0),
    .C(n_3107_o_0),
    .Y(n_3420_o_0));
 OAI311xp33_ASAP7_75t_R n_3421 (.A1(n_3034_o_0),
    .A2(net29),
    .A3(n_3126_o_0),
    .B1(n_3237_o_0),
    .C1(n_3282_o_0),
    .Y(n_3421_o_0));
 OAI221xp5_ASAP7_75t_R n_3422 (.A1(n_3152_o_0),
    .A2(n_3420_o_0),
    .B1(n_3154_o_0),
    .B2(n_3421_o_0),
    .C(n_3269_o_0),
    .Y(n_3422_o_0));
 OAI21xp33_ASAP7_75t_R n_3423 (.A1(n_3417_o_0),
    .A2(n_3419_o_0),
    .B(n_3422_o_0),
    .Y(n_3423_o_0));
 NOR2xp33_ASAP7_75t_R n_3424 (.A(n_3319_o_0),
    .B(n_3104_o_0),
    .Y(n_3424_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3425 (.A1(n_3202_o_0),
    .A2(n_3175_o_0),
    .B(n_3424_o_0),
    .C(n_3154_o_0),
    .Y(n_3425_o_0));
 NAND2xp33_ASAP7_75t_R n_3426 (.A(n_3106_o_0),
    .B(n_3227_o_0),
    .Y(n_3426_o_0));
 AOI21xp33_ASAP7_75t_R n_3427 (.A1(net36),
    .A2(n_3059_o_0),
    .B(n_3124_o_0),
    .Y(n_3427_o_0));
 OAI22xp33_ASAP7_75t_R n_3428 (.A1(n_3426_o_0),
    .A2(n_3232_o_0),
    .B1(n_3147_o_0),
    .B2(n_3427_o_0),
    .Y(n_3428_o_0));
 AOI21xp33_ASAP7_75t_R n_3429 (.A1(n_3122_o_0),
    .A2(n_3428_o_0),
    .B(n_3257_o_0),
    .Y(n_3429_o_0));
 OAI21xp33_ASAP7_75t_R n_3430 (.A1(n_3124_o_0),
    .A2(n_3125_o_0),
    .B(n_3103_o_0),
    .Y(n_3430_o_0));
 AOI21xp33_ASAP7_75t_R n_3431 (.A1(n_3034_o_0),
    .A2(n_3430_o_0),
    .B(n_3245_o_0),
    .Y(n_3431_o_0));
 OAI21xp33_ASAP7_75t_R n_3432 (.A1(n_3131_o_0),
    .A2(net36),
    .B(n_3431_o_0),
    .Y(n_3432_o_0));
 NAND2xp33_ASAP7_75t_R n_3433 (.A(n_3163_o_0),
    .B(n_3107_o_0),
    .Y(n_3433_o_0));
 AOI211xp5_ASAP7_75t_R n_3434 (.A1(n_3433_o_0),
    .A2(n_3132_o_0),
    .B(n_3133_o_0),
    .C(n_3183_o_0),
    .Y(n_3434_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3435 (.A1(n_3010_o_0),
    .A2(n_3133_o_0),
    .B(n_3432_o_0),
    .C(n_3434_o_0),
    .Y(n_3435_o_0));
 AOI211xp5_ASAP7_75t_R n_3436 (.A1(n_3425_o_0),
    .A2(n_3429_o_0),
    .B(n_3435_o_0),
    .C(n_3142_o_0),
    .Y(n_3436_o_0));
 AOI21xp33_ASAP7_75t_R n_3437 (.A1(n_3161_o_0),
    .A2(n_3423_o_0),
    .B(n_3436_o_0),
    .Y(n_3437_o_0));
 OAI211xp5_ASAP7_75t_R n_3438 (.A1(n_3198_o_0),
    .A2(net29),
    .B(n_3184_o_0),
    .C(n_3034_o_0),
    .Y(n_3438_o_0));
 OAI211xp5_ASAP7_75t_R n_3439 (.A1(n_3232_o_0),
    .A2(n_3426_o_0),
    .B(n_3438_o_0),
    .C(n_3133_o_0),
    .Y(n_3439_o_0));
 INVx1_ASAP7_75t_R n_3440 (.A(n_3130_o_0),
    .Y(n_3440_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3441 (.A1(n_3252_o_0),
    .A2(n_3440_o_0),
    .B(n_3178_o_0),
    .C(n_3154_o_0),
    .Y(n_3441_o_0));
 NAND3xp33_ASAP7_75t_R n_3442 (.A(n_3227_o_0),
    .B(n_3430_o_0),
    .C(n_3034_o_0),
    .Y(n_3442_o_0));
 OAI21xp33_ASAP7_75t_R n_3443 (.A1(n_3253_o_0),
    .A2(n_3197_o_0),
    .B(n_3442_o_0),
    .Y(n_3443_o_0));
 OAI31xp33_ASAP7_75t_R n_3444 (.A1(net29),
    .A2(n_3095_o_0),
    .A3(n_3106_o_0),
    .B(n_3151_o_0),
    .Y(n_3444_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3445 (.A1(n_3147_o_0),
    .A2(n_3274_o_0),
    .B(n_3444_o_0),
    .C(n_3269_o_0),
    .Y(n_3445_o_0));
 AOI21xp33_ASAP7_75t_R n_3446 (.A1(n_3122_o_0),
    .A2(n_3443_o_0),
    .B(n_3445_o_0),
    .Y(n_3446_o_0));
 AOI31xp33_ASAP7_75t_R n_3447 (.A1(n_3245_o_0),
    .A2(n_3439_o_0),
    .A3(n_3441_o_0),
    .B(n_3446_o_0),
    .Y(n_3447_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3448 (.A1(n_3147_o_0),
    .A2(n_3164_o_0),
    .B(n_3273_o_0),
    .C(n_3154_o_0),
    .Y(n_3448_o_0));
 AOI311xp33_ASAP7_75t_R n_3449 (.A1(n_3248_o_0),
    .A2(n_3308_o_0),
    .A3(n_3154_o_0),
    .B(n_3234_o_0),
    .C(n_3448_o_0),
    .Y(n_3449_o_0));
 NAND3xp33_ASAP7_75t_R n_3450 (.A(n_3131_o_0),
    .B(n_3106_o_0),
    .C(net29),
    .Y(n_3450_o_0));
 OAI211xp5_ASAP7_75t_R n_3451 (.A1(n_3034_o_0),
    .A2(n_3225_o_0),
    .B(n_3250_o_0),
    .C(n_3450_o_0),
    .Y(n_3451_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3452 (.A1(n_3125_o_0),
    .A2(n_3106_o_0),
    .B(net36),
    .C(n_3151_o_0),
    .Y(n_3452_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3453 (.A1(n_3147_o_0),
    .A2(n_3342_o_0),
    .B(n_3452_o_0),
    .C(n_3245_o_0),
    .Y(n_3453_o_0));
 AOI21xp33_ASAP7_75t_R n_3454 (.A1(n_3133_o_0),
    .A2(n_3451_o_0),
    .B(n_3453_o_0),
    .Y(n_3454_o_0));
 AOI211xp5_ASAP7_75t_R n_3455 (.A1(n_3449_o_0),
    .A2(n_3257_o_0),
    .B(n_3161_o_0),
    .C(n_3454_o_0),
    .Y(n_3455_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3456 (.A1(n_3142_o_0),
    .A2(n_3447_o_0),
    .B(n_3455_o_0),
    .C(n_3020_o_0),
    .Y(n_3456_o_0));
 OAI21xp33_ASAP7_75t_R n_3457 (.A1(n_3020_o_0),
    .A2(n_3437_o_0),
    .B(n_3456_o_0),
    .Y(n_3457_o_0));
 INVx1_ASAP7_75t_R n_3458 (.A(n_3161_o_0),
    .Y(n_3458_o_0));
 OAI21xp33_ASAP7_75t_R n_3459 (.A1(n_3104_o_0),
    .A2(n_3273_o_0),
    .B(n_3282_o_0),
    .Y(n_3459_o_0));
 INVx1_ASAP7_75t_R n_3460 (.A(n_3357_o_0),
    .Y(n_3460_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3461 (.A1(n_3129_o_0),
    .A2(net29),
    .B(n_3290_o_0),
    .C(n_3460_o_0),
    .Y(n_3461_o_0));
 OAI22xp33_ASAP7_75t_R n_3462 (.A1(n_3459_o_0),
    .A2(n_3154_o_0),
    .B1(n_3133_o_0),
    .B2(n_3461_o_0),
    .Y(n_3462_o_0));
 OAI211xp5_ASAP7_75t_R n_3463 (.A1(net36),
    .A2(n_3232_o_0),
    .B(n_3382_o_0),
    .C(n_3107_o_0),
    .Y(n_3463_o_0));
 AOI31xp33_ASAP7_75t_R n_3464 (.A1(n_3106_o_0),
    .A2(n_3259_o_0),
    .A3(n_3189_o_0),
    .B(n_3151_o_0),
    .Y(n_3464_o_0));
 NAND2xp33_ASAP7_75t_R n_3465 (.A(n_3124_o_0),
    .B(n_3034_o_0),
    .Y(n_3465_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3466 (.A1(n_3232_o_0),
    .A2(n_3426_o_0),
    .B(n_3465_o_0),
    .C(n_3133_o_0),
    .Y(n_3466_o_0));
 AOI211xp5_ASAP7_75t_R n_3467 (.A1(n_3463_o_0),
    .A2(n_3464_o_0),
    .B(n_3466_o_0),
    .C(n_3010_o_0),
    .Y(n_3467_o_0));
 AOI21xp33_ASAP7_75t_R n_3468 (.A1(n_3245_o_0),
    .A2(n_3462_o_0),
    .B(n_3467_o_0),
    .Y(n_3468_o_0));
 AOI21xp33_ASAP7_75t_R n_3469 (.A1(net29),
    .A2(n_3126_o_0),
    .B(n_3034_o_0),
    .Y(n_3469_o_0));
 OR3x1_ASAP7_75t_R n_3470 (.A(n_3167_o_0),
    .B(n_3122_o_0),
    .C(n_3395_o_0),
    .Y(n_3470_o_0));
 OAI31xp33_ASAP7_75t_R n_3471 (.A1(n_3154_o_0),
    .A2(n_3254_o_0),
    .A3(n_3469_o_0),
    .B(n_3470_o_0),
    .Y(n_3471_o_0));
 AOI211xp5_ASAP7_75t_R n_3472 (.A1(n_3183_o_0),
    .A2(n_3124_o_0),
    .B(n_3034_o_0),
    .C(n_3111_o_0),
    .Y(n_3472_o_0));
 AOI31xp33_ASAP7_75t_R n_3473 (.A1(n_3034_o_0),
    .A2(n_3125_o_0),
    .A3(n_3218_o_0),
    .B(n_3472_o_0),
    .Y(n_3473_o_0));
 AOI21xp33_ASAP7_75t_R n_3474 (.A1(n_3122_o_0),
    .A2(n_3473_o_0),
    .B(n_3245_o_0),
    .Y(n_3474_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3475 (.A1(n_3127_o_0),
    .A2(n_3185_o_0),
    .B(n_3226_o_0),
    .C(n_3474_o_0),
    .D(n_3142_o_0),
    .Y(n_3475_o_0));
 OAI21xp33_ASAP7_75t_R n_3476 (.A1(n_3257_o_0),
    .A2(n_3471_o_0),
    .B(n_3475_o_0),
    .Y(n_3476_o_0));
 OAI21xp33_ASAP7_75t_R n_3477 (.A1(n_3458_o_0),
    .A2(n_3468_o_0),
    .B(n_3476_o_0),
    .Y(n_3477_o_0));
 OAI21xp33_ASAP7_75t_R n_3478 (.A1(n_3198_o_0),
    .A2(net29),
    .B(n_3290_o_0),
    .Y(n_3478_o_0));
 OA21x2_ASAP7_75t_R n_3479 (.A1(n_3203_o_0),
    .A2(n_3342_o_0),
    .B(n_3478_o_0),
    .Y(n_3479_o_0));
 OAI31xp33_ASAP7_75t_R n_3480 (.A1(n_3185_o_0),
    .A2(n_3236_o_0),
    .A3(n_3245_o_0),
    .B(n_3122_o_0),
    .Y(n_3480_o_0));
 AOI21xp33_ASAP7_75t_R n_3481 (.A1(n_3010_o_0),
    .A2(n_3479_o_0),
    .B(n_3480_o_0),
    .Y(n_3481_o_0));
 INVx1_ASAP7_75t_R n_3482 (.A(n_3266_o_0),
    .Y(n_3482_o_0));
 OAI21xp33_ASAP7_75t_R n_3483 (.A1(n_3147_o_0),
    .A2(n_3168_o_0),
    .B(n_3482_o_0),
    .Y(n_3483_o_0));
 OAI22xp33_ASAP7_75t_R n_3484 (.A1(n_3482_o_0),
    .A2(n_3191_o_0),
    .B1(n_3010_o_0),
    .B2(n_3329_o_0),
    .Y(n_3484_o_0));
 AOI21xp33_ASAP7_75t_R n_3485 (.A1(n_3245_o_0),
    .A2(n_3483_o_0),
    .B(n_3484_o_0),
    .Y(n_3485_o_0));
 OAI21xp33_ASAP7_75t_R n_3486 (.A1(n_3133_o_0),
    .A2(n_3485_o_0),
    .B(n_3142_o_0),
    .Y(n_3486_o_0));
 AOI21xp33_ASAP7_75t_R n_3487 (.A1(n_3394_o_0),
    .A2(n_3266_o_0),
    .B(n_3257_o_0),
    .Y(n_3487_o_0));
 OAI21xp33_ASAP7_75t_R n_3488 (.A1(n_3382_o_0),
    .A2(n_3147_o_0),
    .B(n_3487_o_0),
    .Y(n_3488_o_0));
 AOI31xp33_ASAP7_75t_R n_3489 (.A1(n_3147_o_0),
    .A2(n_3382_o_0),
    .A3(n_3227_o_0),
    .B(n_3245_o_0),
    .Y(n_3489_o_0));
 OAI21xp33_ASAP7_75t_R n_3490 (.A1(n_3239_o_0),
    .A2(n_3191_o_0),
    .B(n_3489_o_0),
    .Y(n_3490_o_0));
 OAI211xp5_ASAP7_75t_R n_3491 (.A1(n_3259_o_0),
    .A2(net36),
    .B(n_3034_o_0),
    .C(n_3189_o_0),
    .Y(n_3491_o_0));
 AOI22xp33_ASAP7_75t_R n_3492 (.A1(n_3301_o_0),
    .A2(n_3210_o_0),
    .B1(n_3145_o_0),
    .B2(n_3059_o_0),
    .Y(n_3492_o_0));
 NAND2xp33_ASAP7_75t_R n_3493 (.A(n_3245_o_0),
    .B(n_3151_o_0),
    .Y(n_3493_o_0));
 NAND2xp33_ASAP7_75t_R n_3494 (.A(n_3059_o_0),
    .B(n_3034_o_0),
    .Y(n_3494_o_0));
 INVx1_ASAP7_75t_R n_3495 (.A(n_3494_o_0),
    .Y(n_3495_o_0));
 NOR2xp33_ASAP7_75t_R n_3496 (.A(n_3010_o_0),
    .B(n_3133_o_0),
    .Y(n_3496_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3497 (.A1(n_3173_o_0),
    .A2(n_3175_o_0),
    .B(n_3495_o_0),
    .C(n_3496_o_0),
    .Y(n_3497_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3498 (.A1(n_3491_o_0),
    .A2(n_3492_o_0),
    .B(n_3493_o_0),
    .C(n_3497_o_0),
    .Y(n_3498_o_0));
 AOI31xp33_ASAP7_75t_R n_3499 (.A1(n_3122_o_0),
    .A2(n_3488_o_0),
    .A3(n_3490_o_0),
    .B(n_3498_o_0),
    .Y(n_3499_o_0));
 AOI21xp33_ASAP7_75t_R n_3500 (.A1(n_3458_o_0),
    .A2(n_3499_o_0),
    .B(n_3241_o_0),
    .Y(n_3500_o_0));
 OAI21xp33_ASAP7_75t_R n_3501 (.A1(n_3481_o_0),
    .A2(n_3486_o_0),
    .B(n_3500_o_0),
    .Y(n_3501_o_0));
 OAI21xp33_ASAP7_75t_R n_3502 (.A1(n_3020_o_0),
    .A2(n_3477_o_0),
    .B(n_3501_o_0),
    .Y(n_3502_o_0));
 NOR2xp33_ASAP7_75t_R n_3503 (.A(n_3133_o_0),
    .B(n_3269_o_0),
    .Y(n_3503_o_0));
 AOI21xp33_ASAP7_75t_R n_3504 (.A1(n_3394_o_0),
    .A2(n_3272_o_0),
    .B(n_3151_o_0),
    .Y(n_3504_o_0));
 OAI31xp33_ASAP7_75t_R n_3505 (.A1(n_3125_o_0),
    .A2(net29),
    .A3(n_3107_o_0),
    .B(n_3504_o_0),
    .Y(n_3505_o_0));
 OAI33xp33_ASAP7_75t_R n_3506 (.A1(net40),
    .A2(n_3102_o_0),
    .A3(n_3110_o_0),
    .B1(n_3076_o_0),
    .B2(n_3103_o_0),
    .B3(n_3162_o_0),
    .Y(n_3506_o_0));
 INVx1_ASAP7_75t_R n_3507 (.A(n_3506_o_0),
    .Y(n_3507_o_0));
 AOI31xp33_ASAP7_75t_R n_3508 (.A1(n_3147_o_0),
    .A2(n_3382_o_0),
    .A3(n_3227_o_0),
    .B(n_3122_o_0),
    .Y(n_3508_o_0));
 OAI21xp33_ASAP7_75t_R n_3509 (.A1(n_3147_o_0),
    .A2(n_3507_o_0),
    .B(n_3508_o_0),
    .Y(n_3509_o_0));
 NAND4xp25_ASAP7_75t_R n_3510 (.A(n_3442_o_0),
    .B(n_3153_o_0),
    .C(n_3133_o_0),
    .D(n_3010_o_0),
    .Y(n_3510_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3511 (.A1(n_3505_o_0),
    .A2(n_3509_o_0),
    .B(n_3245_o_0),
    .C(n_3510_o_0),
    .Y(n_3511_o_0));
 AOI21xp33_ASAP7_75t_R n_3512 (.A1(n_3345_o_0),
    .A2(n_3503_o_0),
    .B(n_3511_o_0),
    .Y(n_3512_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3513 (.A1(n_3107_o_0),
    .A2(n_3275_o_0),
    .B(n_3319_o_0),
    .C(n_3214_o_0),
    .Y(n_3513_o_0));
 AOI21xp33_ASAP7_75t_R n_3514 (.A1(net40),
    .A2(n_3494_o_0),
    .B(n_3122_o_0),
    .Y(n_3514_o_0));
 OAI21xp33_ASAP7_75t_R n_3515 (.A1(n_3125_o_0),
    .A2(net29),
    .B(n_3514_o_0),
    .Y(n_3515_o_0));
 OAI21xp33_ASAP7_75t_R n_3516 (.A1(n_3151_o_0),
    .A2(n_3513_o_0),
    .B(n_3515_o_0),
    .Y(n_3516_o_0));
 OAI211xp5_ASAP7_75t_R n_3517 (.A1(n_3183_o_0),
    .A2(n_3181_o_0),
    .B(n_3433_o_0),
    .C(n_3133_o_0),
    .Y(n_3517_o_0));
 AOI211xp5_ASAP7_75t_R n_3518 (.A1(n_3281_o_0),
    .A2(n_3145_o_0),
    .B(n_3395_o_0),
    .C(n_3133_o_0),
    .Y(n_3518_o_0));
 INVx1_ASAP7_75t_R n_3519 (.A(n_3518_o_0),
    .Y(n_3519_o_0));
 AOI21xp33_ASAP7_75t_R n_3520 (.A1(n_3517_o_0),
    .A2(n_3519_o_0),
    .B(n_3269_o_0),
    .Y(n_3520_o_0));
 AOI211xp5_ASAP7_75t_R n_3521 (.A1(n_3269_o_0),
    .A2(n_3516_o_0),
    .B(n_3520_o_0),
    .C(n_3142_o_0),
    .Y(n_3521_o_0));
 AOI21xp33_ASAP7_75t_R n_3522 (.A1(n_3161_o_0),
    .A2(n_3512_o_0),
    .B(n_3521_o_0),
    .Y(n_3522_o_0));
 AO21x1_ASAP7_75t_R n_3523 (.A1(n_3147_o_0),
    .A2(n_3166_o_0),
    .B(n_3010_o_0),
    .Y(n_3523_o_0));
 INVx1_ASAP7_75t_R n_3524 (.A(n_3334_o_0),
    .Y(n_3524_o_0));
 OAI211xp5_ASAP7_75t_R n_3525 (.A1(n_3059_o_0),
    .A2(net40),
    .B(n_3107_o_0),
    .C(n_3163_o_0),
    .Y(n_3525_o_0));
 OAI31xp33_ASAP7_75t_R n_3526 (.A1(n_3168_o_0),
    .A2(n_3107_o_0),
    .A3(net29),
    .B(n_3525_o_0),
    .Y(n_3526_o_0));
 AOI21xp33_ASAP7_75t_R n_3527 (.A1(n_3245_o_0),
    .A2(n_3526_o_0),
    .B(n_3151_o_0),
    .Y(n_3527_o_0));
 OAI21xp33_ASAP7_75t_R n_3528 (.A1(n_3523_o_0),
    .A2(n_3524_o_0),
    .B(n_3527_o_0),
    .Y(n_3528_o_0));
 OAI21xp33_ASAP7_75t_R n_3529 (.A1(n_3248_o_0),
    .A2(n_3129_o_0),
    .B(n_3308_o_0),
    .Y(n_3529_o_0));
 OAI31xp33_ASAP7_75t_R n_3530 (.A1(n_3147_o_0),
    .A2(n_3148_o_0),
    .A3(n_3176_o_0),
    .B(n_3529_o_0),
    .Y(n_3530_o_0));
 INVx1_ASAP7_75t_R n_3531 (.A(n_3530_o_0),
    .Y(n_3531_o_0));
 AO21x1_ASAP7_75t_R n_3532 (.A1(n_3131_o_0),
    .A2(net36),
    .B(n_3203_o_0),
    .Y(n_3532_o_0));
 OAI31xp33_ASAP7_75t_R n_3533 (.A1(n_3147_o_0),
    .A2(n_3191_o_0),
    .A3(n_3228_o_0),
    .B(n_3532_o_0),
    .Y(n_3533_o_0));
 AOI21xp33_ASAP7_75t_R n_3534 (.A1(n_3257_o_0),
    .A2(n_3533_o_0),
    .B(n_3133_o_0),
    .Y(n_3534_o_0));
 OAI21xp33_ASAP7_75t_R n_3535 (.A1(n_3257_o_0),
    .A2(n_3531_o_0),
    .B(n_3534_o_0),
    .Y(n_3535_o_0));
 AOI31xp33_ASAP7_75t_R n_3536 (.A1(n_3528_o_0),
    .A2(n_3535_o_0),
    .A3(n_3142_o_0),
    .B(n_3020_o_0),
    .Y(n_3536_o_0));
 AOI21xp33_ASAP7_75t_R n_3537 (.A1(n_3106_o_0),
    .A2(n_3280_o_0),
    .B(n_3356_o_0),
    .Y(n_3537_o_0));
 AOI211xp5_ASAP7_75t_R n_3538 (.A1(n_3107_o_0),
    .A2(n_3268_o_0),
    .B(n_3537_o_0),
    .C(n_3010_o_0),
    .Y(n_3538_o_0));
 NOR2xp33_ASAP7_75t_R n_3539 (.A(n_3010_o_0),
    .B(n_3133_o_0),
    .Y(n_3539_o_0));
 INVx1_ASAP7_75t_R n_3540 (.A(n_3177_o_0),
    .Y(n_3540_o_0));
 AOI22xp33_ASAP7_75t_R n_3541 (.A1(n_3540_o_0),
    .A2(n_3249_o_0),
    .B1(n_3147_o_0),
    .B2(net40),
    .Y(n_3541_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3542 (.A1(n_3133_o_0),
    .A2(n_3538_o_0),
    .B(n_3539_o_0),
    .C(n_3541_o_0),
    .D(n_3122_o_0),
    .Y(n_3542_o_0));
 AOI211xp5_ASAP7_75t_R n_3543 (.A1(n_3538_o_0),
    .A2(n_3133_o_0),
    .B(n_3154_o_0),
    .C(n_3539_o_0),
    .Y(n_3543_o_0));
 NOR3xp33_ASAP7_75t_R n_3544 (.A(n_3275_o_0),
    .B(n_3387_o_0),
    .C(n_3107_o_0),
    .Y(n_3544_o_0));
 AOI31xp33_ASAP7_75t_R n_3545 (.A1(n_3034_o_0),
    .A2(n_3440_o_0),
    .A3(n_3165_o_0),
    .B(n_3544_o_0),
    .Y(n_3545_o_0));
 NOR3xp33_ASAP7_75t_R n_3546 (.A(n_3095_o_0),
    .B(net29),
    .C(n_3034_o_0),
    .Y(n_3546_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3547 (.A1(net29),
    .A2(n_3059_o_0),
    .B(n_3356_o_0),
    .C(n_3546_o_0),
    .Y(n_3547_o_0));
 NAND2xp33_ASAP7_75t_R n_3548 (.A(n_3059_o_0),
    .B(n_3145_o_0),
    .Y(n_3548_o_0));
 AOI31xp33_ASAP7_75t_R n_3549 (.A1(n_3122_o_0),
    .A2(n_3547_o_0),
    .A3(n_3548_o_0),
    .B(n_3257_o_0),
    .Y(n_3549_o_0));
 OAI21xp33_ASAP7_75t_R n_3550 (.A1(n_3133_o_0),
    .A2(n_3545_o_0),
    .B(n_3549_o_0),
    .Y(n_3550_o_0));
 OAI211xp5_ASAP7_75t_R n_3551 (.A1(n_3542_o_0),
    .A2(n_3543_o_0),
    .B(n_3550_o_0),
    .C(n_3143_o_0),
    .Y(n_3551_o_0));
 AOI22xp33_ASAP7_75t_R n_3552 (.A1(n_3522_o_0),
    .A2(n_3020_o_0),
    .B1(n_3536_o_0),
    .B2(n_3551_o_0),
    .Y(n_3552_o_0));
 AOI31xp33_ASAP7_75t_R n_3553 (.A1(n_3034_o_0),
    .A2(n_3184_o_0),
    .A3(n_3225_o_0),
    .B(n_3544_o_0),
    .Y(n_3553_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3554 (.A1(n_3107_o_0),
    .A2(n_3275_o_0),
    .B(n_3442_o_0),
    .C(n_3010_o_0),
    .Y(n_3554_o_0));
 INVx1_ASAP7_75t_R n_3555 (.A(n_3554_o_0),
    .Y(n_3555_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3556 (.A1(n_3269_o_0),
    .A2(n_3553_o_0),
    .B(n_3555_o_0),
    .C(n_3133_o_0),
    .Y(n_3556_o_0));
 OAI32xp33_ASAP7_75t_R n_3557 (.A1(n_3147_o_0),
    .A2(n_3297_o_0),
    .A3(n_3275_o_0),
    .B1(n_3190_o_0),
    .B2(n_3166_o_0),
    .Y(n_3557_o_0));
 INVx1_ASAP7_75t_R n_3558 (.A(n_3557_o_0),
    .Y(n_3558_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3559 (.A1(n_3125_o_0),
    .A2(net40),
    .B(net36),
    .C(n_3215_o_0),
    .Y(n_3559_o_0));
 INVx1_ASAP7_75t_R n_3560 (.A(n_3559_o_0),
    .Y(n_3560_o_0));
 OAI21xp33_ASAP7_75t_R n_3561 (.A1(n_3148_o_0),
    .A2(n_3190_o_0),
    .B(n_3269_o_0),
    .Y(n_3561_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3562 (.A1(n_3560_o_0),
    .A2(n_3107_o_0),
    .B(n_3561_o_0),
    .C(n_3133_o_0),
    .Y(n_3562_o_0));
 AOI21xp33_ASAP7_75t_R n_3563 (.A1(n_3245_o_0),
    .A2(n_3558_o_0),
    .B(n_3562_o_0),
    .Y(n_3563_o_0));
 NOR2xp33_ASAP7_75t_R n_3564 (.A(n_3319_o_0),
    .B(n_3104_o_0),
    .Y(n_3564_o_0));
 AOI311xp33_ASAP7_75t_R n_3565 (.A1(n_3106_o_0),
    .A2(n_3165_o_0),
    .A3(n_3227_o_0),
    .B(n_3245_o_0),
    .C(n_3564_o_0),
    .Y(n_3565_o_0));
 AOI211xp5_ASAP7_75t_R n_3566 (.A1(n_3147_o_0),
    .A2(n_3166_o_0),
    .B(n_3255_o_0),
    .C(n_3269_o_0),
    .Y(n_3566_o_0));
 OAI22xp33_ASAP7_75t_R n_3567 (.A1(n_3164_o_0),
    .A2(n_3203_o_0),
    .B1(n_3147_o_0),
    .B2(n_3148_o_0),
    .Y(n_3567_o_0));
 INVx1_ASAP7_75t_R n_3568 (.A(n_3163_o_0),
    .Y(n_3568_o_0));
 OAI31xp33_ASAP7_75t_R n_3569 (.A1(n_3106_o_0),
    .A2(n_3568_o_0),
    .A3(n_3183_o_0),
    .B(n_3269_o_0),
    .Y(n_3569_o_0));
 AOI21xp33_ASAP7_75t_R n_3570 (.A1(n_3125_o_0),
    .A2(n_3106_o_0),
    .B(n_3569_o_0),
    .Y(n_3570_o_0));
 AOI21xp33_ASAP7_75t_R n_3571 (.A1(n_3010_o_0),
    .A2(n_3567_o_0),
    .B(n_3570_o_0),
    .Y(n_3571_o_0));
 OAI321xp33_ASAP7_75t_R n_3572 (.A1(n_3565_o_0),
    .A2(n_3566_o_0),
    .A3(n_3122_o_0),
    .B1(n_3571_o_0),
    .B2(n_3151_o_0),
    .C(n_3161_o_0),
    .Y(n_3572_o_0));
 OAI31xp33_ASAP7_75t_R n_3573 (.A1(n_3142_o_0),
    .A2(n_3556_o_0),
    .A3(n_3563_o_0),
    .B(n_3572_o_0),
    .Y(n_3573_o_0));
 AOI21xp33_ASAP7_75t_R n_3574 (.A1(n_3237_o_0),
    .A2(n_3296_o_0),
    .B(n_3034_o_0),
    .Y(n_3574_o_0));
 AOI31xp33_ASAP7_75t_R n_3575 (.A1(net40),
    .A2(net36),
    .A3(n_3107_o_0),
    .B(n_3574_o_0),
    .Y(n_3575_o_0));
 AOI21xp33_ASAP7_75t_R n_3576 (.A1(n_3059_o_0),
    .A2(n_3163_o_0),
    .B(net40),
    .Y(n_3576_o_0));
 OAI211xp5_ASAP7_75t_R n_3577 (.A1(n_3034_o_0),
    .A2(n_3576_o_0),
    .B(n_3250_o_0),
    .C(n_3122_o_0),
    .Y(n_3577_o_0));
 OAI21xp33_ASAP7_75t_R n_3578 (.A1(n_3274_o_0),
    .A2(n_3106_o_0),
    .B(n_3217_o_0),
    .Y(n_3578_o_0));
 INVx1_ASAP7_75t_R n_3579 (.A(n_3189_o_0),
    .Y(n_3579_o_0));
 NAND2xp33_ASAP7_75t_R n_3580 (.A(n_3296_o_0),
    .B(n_3272_o_0),
    .Y(n_3580_o_0));
 OAI31xp33_ASAP7_75t_R n_3581 (.A1(n_3107_o_0),
    .A2(n_3579_o_0),
    .A3(n_3228_o_0),
    .B(n_3580_o_0),
    .Y(n_3581_o_0));
 NOR2xp33_ASAP7_75t_R n_3582 (.A(n_3154_o_0),
    .B(n_3269_o_0),
    .Y(n_3582_o_0));
 AOI321xp33_ASAP7_75t_R n_3583 (.A1(n_3269_o_0),
    .A2(n_3577_o_0),
    .A3(n_3578_o_0),
    .B1(n_3581_o_0),
    .B2(n_3582_o_0),
    .C(n_3143_o_0),
    .Y(n_3583_o_0));
 OAI31xp33_ASAP7_75t_R n_3584 (.A1(n_3575_o_0),
    .A2(n_3269_o_0),
    .A3(n_3133_o_0),
    .B(n_3583_o_0),
    .Y(n_3584_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3585 (.A1(net29),
    .A2(n_3198_o_0),
    .B(n_3272_o_0),
    .C(n_3133_o_0),
    .Y(n_3585_o_0));
 OA21x2_ASAP7_75t_R n_3586 (.A1(n_3034_o_0),
    .A2(n_3559_o_0),
    .B(n_3585_o_0),
    .Y(n_3586_o_0));
 NOR2xp33_ASAP7_75t_R n_3587 (.A(n_3387_o_0),
    .B(n_3329_o_0),
    .Y(n_3587_o_0));
 AOI31xp33_ASAP7_75t_R n_3588 (.A1(n_3106_o_0),
    .A2(n_3287_o_0),
    .A3(n_3259_o_0),
    .B(n_3587_o_0),
    .Y(n_3588_o_0));
 AO21x1_ASAP7_75t_R n_3589 (.A1(n_3588_o_0),
    .A2(n_3133_o_0),
    .B(n_3010_o_0),
    .Y(n_3589_o_0));
 OAI211xp5_ASAP7_75t_R n_3590 (.A1(n_3106_o_0),
    .A2(n_3225_o_0),
    .B(n_3217_o_0),
    .C(n_3280_o_0),
    .Y(n_3590_o_0));
 AOI21xp33_ASAP7_75t_R n_3591 (.A1(n_3147_o_0),
    .A2(n_3301_o_0),
    .B(n_3154_o_0),
    .Y(n_3591_o_0));
 OAI21xp33_ASAP7_75t_R n_3592 (.A1(n_3380_o_0),
    .A2(n_3177_o_0),
    .B(n_3591_o_0),
    .Y(n_3592_o_0));
 AOI31xp33_ASAP7_75t_R n_3593 (.A1(n_3010_o_0),
    .A2(n_3590_o_0),
    .A3(n_3592_o_0),
    .B(n_3142_o_0),
    .Y(n_3593_o_0));
 OAI21xp33_ASAP7_75t_R n_3594 (.A1(n_3586_o_0),
    .A2(n_3589_o_0),
    .B(n_3593_o_0),
    .Y(n_3594_o_0));
 OAI211xp5_ASAP7_75t_R n_3595 (.A1(n_3017_o_0),
    .A2(n_3019_o_0),
    .B(n_3584_o_0),
    .C(n_3594_o_0),
    .Y(n_3595_o_0));
 OAI21xp33_ASAP7_75t_R n_3596 (.A1(n_3241_o_0),
    .A2(n_3573_o_0),
    .B(n_3595_o_0),
    .Y(n_3596_o_0));
 XNOR2xp5_ASAP7_75t_R n_3597 (.A(_01008_),
    .B(_01048_),
    .Y(n_3597_o_0));
 XNOR2xp5_ASAP7_75t_R n_3598 (.A(_01088_),
    .B(_01096_),
    .Y(n_3598_o_0));
 XNOR2xp5_ASAP7_75t_R n_3599 (.A(_01049_),
    .B(n_3598_o_0),
    .Y(n_3599_o_0));
 XOR2xp5_ASAP7_75t_R n_3600 (.A(n_3597_o_0),
    .B(n_3599_o_0),
    .Y(n_3600_o_0));
 NOR2xp33_ASAP7_75t_R n_3601 (.A(_00671_),
    .B(net),
    .Y(n_3601_o_0));
 AOI21xp33_ASAP7_75t_R n_3602 (.A1(net),
    .A2(n_3600_o_0),
    .B(n_3601_o_0),
    .Y(n_3602_o_0));
 NAND2xp33_ASAP7_75t_R n_3603 (.A(_00921_),
    .B(n_3602_o_0),
    .Y(n_3603_o_0));
 OAI21xp33_ASAP7_75t_R n_3604 (.A1(_00921_),
    .A2(n_3602_o_0),
    .B(n_3603_o_0),
    .Y(n_3604_o_0));
 INVx1_ASAP7_75t_R n_3605 (.A(n_3604_o_0),
    .Y(n_3605_o_0));
 XOR2xp5_ASAP7_75t_R n_3606 (.A(_01010_),
    .B(_01050_),
    .Y(n_3606_o_0));
 XNOR2xp5_ASAP7_75t_R n_3607 (.A(_01051_),
    .B(_01090_),
    .Y(n_3607_o_0));
 XNOR2xp5_ASAP7_75t_R n_3608 (.A(_01098_),
    .B(n_3607_o_0),
    .Y(n_3608_o_0));
 NOR2xp33_ASAP7_75t_R n_3609 (.A(n_3606_o_0),
    .B(n_3608_o_0),
    .Y(n_3609_o_0));
 NOR2xp33_ASAP7_75t_R n_3610 (.A(_00669_),
    .B(net),
    .Y(n_3610_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3611 (.A1(n_3606_o_0),
    .A2(n_3608_o_0),
    .B(n_3609_o_0),
    .C(net),
    .D(n_3610_o_0),
    .Y(n_3611_o_0));
 NAND2xp33_ASAP7_75t_R n_3612 (.A(_00923_),
    .B(n_3611_o_0),
    .Y(n_3612_o_0));
 OAI21xp33_ASAP7_75t_R n_3613 (.A1(_00923_),
    .A2(n_3611_o_0),
    .B(n_3612_o_0),
    .Y(n_3613_o_0));
 XOR2xp5_ASAP7_75t_R n_3614 (.A(_01006_),
    .B(_01011_),
    .Y(n_3614_o_0));
 XNOR2xp5_ASAP7_75t_R n_3615 (.A(_01047_),
    .B(n_3614_o_0),
    .Y(n_3615_o_0));
 XNOR2xp5_ASAP7_75t_R n_3616 (.A(_01046_),
    .B(_01051_),
    .Y(n_3616_o_0));
 XNOR2xp5_ASAP7_75t_R n_3617 (.A(_01086_),
    .B(_01094_),
    .Y(n_3617_o_0));
 XNOR2xp5_ASAP7_75t_R n_3618 (.A(n_3616_o_0),
    .B(n_3617_o_0),
    .Y(n_3618_o_0));
 NAND2xp33_ASAP7_75t_R n_3619 (.A(n_3618_o_0),
    .B(n_3615_o_0),
    .Y(n_3619_o_0));
 OAI21xp33_ASAP7_75t_R n_3620 (.A1(n_3615_o_0),
    .A2(n_3618_o_0),
    .B(n_3619_o_0),
    .Y(n_3620_o_0));
 NOR2xp33_ASAP7_75t_R n_3621 (.A(_00673_),
    .B(net77),
    .Y(n_3621_o_0));
 AOI211xp5_ASAP7_75t_R n_3622 (.A1(n_3620_o_0),
    .A2(net77),
    .B(_00919_),
    .C(n_3621_o_0),
    .Y(n_3622_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3623 (.A1(n_3620_o_0),
    .A2(net39),
    .B(n_3621_o_0),
    .C(_00919_),
    .D(n_3622_o_0),
    .Y(n_3623_o_0));
 INVx2_ASAP7_75t_R n_3624 (.A(n_3623_o_0),
    .Y(n_3624_o_0));
 AOI211xp5_ASAP7_75t_R n_3625 (.A1(n_3620_o_0),
    .A2(net39),
    .B(n_2399_o_0),
    .C(n_3621_o_0),
    .Y(n_3625_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3626 (.A1(net39),
    .A2(n_3620_o_0),
    .B(n_3621_o_0),
    .C(n_2399_o_0),
    .D(n_3625_o_0),
    .Y(n_3626_o_0));
 INVx3_ASAP7_75t_R n_3627 (.A(n_3626_o_0),
    .Y(n_3627_o_0));
 INVx1_ASAP7_75t_R n_3628 (.A(_00502_),
    .Y(n_3628_o_0));
 XNOR2xp5_ASAP7_75t_R n_3629 (.A(_01005_),
    .B(_01045_),
    .Y(n_3629_o_0));
 INVx1_ASAP7_75t_R n_3630 (.A(n_3629_o_0),
    .Y(n_3630_o_0));
 XNOR2xp5_ASAP7_75t_R n_3631 (.A(_01085_),
    .B(_01093_),
    .Y(n_3631_o_0));
 XNOR2xp5_ASAP7_75t_R n_3632 (.A(_01046_),
    .B(n_3631_o_0),
    .Y(n_3632_o_0));
 NAND2xp33_ASAP7_75t_R n_3633 (.A(n_3630_o_0),
    .B(n_3632_o_0),
    .Y(n_3633_o_0));
 XOR2xp5_ASAP7_75t_R n_3634 (.A(_01046_),
    .B(n_3631_o_0),
    .Y(n_3634_o_0));
 AOI21xp33_ASAP7_75t_R n_3635 (.A1(n_3629_o_0),
    .A2(n_3634_o_0),
    .B(net3),
    .Y(n_3635_o_0));
 AOI21xp33_ASAP7_75t_R n_3636 (.A1(n_3633_o_0),
    .A2(n_3635_o_0),
    .B(n_2463_o_0),
    .Y(n_3636_o_0));
 OAI21xp33_ASAP7_75t_R n_3637 (.A1(n_3628_o_0),
    .A2(net39),
    .B(n_3636_o_0),
    .Y(n_3637_o_0));
 XNOR2xp5_ASAP7_75t_R n_3638 (.A(n_3629_o_0),
    .B(n_3632_o_0),
    .Y(n_3638_o_0));
 OAI21xp33_ASAP7_75t_R n_3639 (.A1(_00502_),
    .A2(net39),
    .B(n_2463_o_0),
    .Y(n_3639_o_0));
 INVx1_ASAP7_75t_R n_3640 (.A(n_3639_o_0),
    .Y(n_3640_o_0));
 OAI21xp33_ASAP7_75t_R n_3641 (.A1(net5),
    .A2(n_3638_o_0),
    .B(n_3640_o_0),
    .Y(n_3641_o_0));
 NAND2xp5_ASAP7_75t_R n_3642 (.A(n_3637_o_0),
    .B(n_3641_o_0),
    .Y(n_3642_o_0));
 XNOR2xp5_ASAP7_75t_R n_3643 (.A(_01004_),
    .B(_01011_),
    .Y(n_3643_o_0));
 NAND2xp33_ASAP7_75t_R n_3644 (.A(_01092_),
    .B(n_3643_o_0),
    .Y(n_3644_o_0));
 OA21x2_ASAP7_75t_R n_3645 (.A1(_01092_),
    .A2(n_3643_o_0),
    .B(n_3644_o_0),
    .Y(n_3645_o_0));
 XNOR2xp5_ASAP7_75t_R n_3646 (.A(_01045_),
    .B(_01084_),
    .Y(n_3646_o_0));
 XNOR2xp5_ASAP7_75t_R n_3647 (.A(_01044_),
    .B(_01051_),
    .Y(n_3647_o_0));
 XOR2xp5_ASAP7_75t_R n_3648 (.A(n_3646_o_0),
    .B(n_3647_o_0),
    .Y(n_3648_o_0));
 OAI211xp5_ASAP7_75t_R n_3649 (.A1(_01092_),
    .A2(n_3643_o_0),
    .B(n_3648_o_0),
    .C(n_3644_o_0),
    .Y(n_3649_o_0));
 OAI21xp33_ASAP7_75t_R n_3650 (.A1(n_3645_o_0),
    .A2(n_3648_o_0),
    .B(n_3649_o_0),
    .Y(n_3650_o_0));
 OAI21xp33_ASAP7_75t_R n_3651 (.A1(_00499_),
    .A2(net39),
    .B(_00917_),
    .Y(n_3651_o_0));
 INVx1_ASAP7_75t_R n_3652 (.A(n_3651_o_0),
    .Y(n_3652_o_0));
 INVx1_ASAP7_75t_R n_3653 (.A(_01004_),
    .Y(n_3653_o_0));
 NAND2xp33_ASAP7_75t_R n_3654 (.A(_01011_),
    .B(n_3653_o_0),
    .Y(n_3654_o_0));
 OR2x2_ASAP7_75t_R n_3655 (.A(_01011_),
    .B(n_3653_o_0),
    .Y(n_3655_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3656 (.A1(n_3654_o_0),
    .A2(n_3655_o_0),
    .B(_01092_),
    .C(n_3644_o_0),
    .D(n_3648_o_0),
    .Y(n_3656_o_0));
 AO21x1_ASAP7_75t_R n_3657 (.A1(n_3021_o_0),
    .A2(_00499_),
    .B(_00917_),
    .Y(n_3657_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3658 (.A1(n_3645_o_0),
    .A2(n_3648_o_0),
    .B(n_3656_o_0),
    .C(net39),
    .D(n_3657_o_0),
    .Y(n_3658_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_3659 (.A1(n_3021_o_0),
    .A2(n_3650_o_0),
    .B(n_3652_o_0),
    .C(n_3658_o_0),
    .Y(n_3659_o_0));
 INVx1_ASAP7_75t_R n_3660 (.A(n_3659_o_0),
    .Y(n_3660_o_0));
 NAND2xp33_ASAP7_75t_R n_3661 (.A(n_3642_o_0),
    .B(n_3660_o_0),
    .Y(n_3661_o_0));
 NAND2xp33_ASAP7_75t_R n_3662 (.A(n_3627_o_0),
    .B(n_3661_o_0),
    .Y(n_3662_o_0));
 INVx1_ASAP7_75t_R n_3663 (.A(_01091_),
    .Y(n_3663_o_0));
 XNOR2xp5_ASAP7_75t_R n_3664 (.A(_01011_),
    .B(_01051_),
    .Y(n_3664_o_0));
 OR2x2_ASAP7_75t_R n_3665 (.A(n_3663_o_0),
    .B(n_3664_o_0),
    .Y(n_3665_o_0));
 NAND2xp33_ASAP7_75t_R n_3666 (.A(n_3663_o_0),
    .B(n_3664_o_0),
    .Y(n_3666_o_0));
 XNOR2xp5_ASAP7_75t_R n_3667 (.A(_01044_),
    .B(_01083_),
    .Y(n_3667_o_0));
 INVx1_ASAP7_75t_R n_3668 (.A(n_3667_o_0),
    .Y(n_3668_o_0));
 OAI211xp5_ASAP7_75t_R n_3669 (.A1(n_3664_o_0),
    .A2(n_3663_o_0),
    .B(n_3666_o_0),
    .C(n_3668_o_0),
    .Y(n_3669_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3670 (.A1(n_3665_o_0),
    .A2(n_3666_o_0),
    .B(n_3668_o_0),
    .C(n_3669_o_0),
    .Y(n_3670_o_0));
 NOR2xp33_ASAP7_75t_R n_3671 (.A(_00500_),
    .B(net77),
    .Y(n_3671_o_0));
 AOI211xp5_ASAP7_75t_R n_3672 (.A1(n_3670_o_0),
    .A2(net77),
    .B(n_2421_o_0),
    .C(n_3671_o_0),
    .Y(n_3672_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3673 (.A1(net39),
    .A2(n_3670_o_0),
    .B(n_3671_o_0),
    .C(n_2421_o_0),
    .D(n_3672_o_0),
    .Y(n_3673_o_0));
 AOI21xp33_ASAP7_75t_R n_3674 (.A1(n_3628_o_0),
    .A2(net2),
    .B(_00918_),
    .Y(n_3674_o_0));
 AOI221xp5_ASAP7_75t_R n_3675 (.A1(_00502_),
    .A2(net2),
    .B1(n_3633_o_0),
    .B2(n_3635_o_0),
    .C(n_2463_o_0),
    .Y(n_3675_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3676 (.A1(n_3638_o_0),
    .A2(net2),
    .B(n_3674_o_0),
    .C(n_3675_o_0),
    .Y(n_3676_o_0));
 OAI21xp33_ASAP7_75t_R n_3677 (.A1(net2),
    .A2(n_3650_o_0),
    .B(n_3652_o_0),
    .Y(n_3677_o_0));
 INVx1_ASAP7_75t_R n_3678 (.A(n_3658_o_0),
    .Y(n_3678_o_0));
 NAND3xp33_ASAP7_75t_R n_3679 (.A(n_3676_o_0),
    .B(n_3677_o_0),
    .C(n_3678_o_0),
    .Y(n_3679_o_0));
 NOR2xp33_ASAP7_75t_R n_3680 (.A(net50),
    .B(n_3679_o_0),
    .Y(n_3680_o_0));
 NOR2xp33_ASAP7_75t_R n_3681 (.A(n_3630_o_0),
    .B(n_3632_o_0),
    .Y(n_3681_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3682 (.A1(n_3630_o_0),
    .A2(n_3632_o_0),
    .B(n_3681_o_0),
    .C(net77),
    .D(n_3639_o_0),
    .Y(n_3682_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_3683 (.A1(n_3628_o_0),
    .A2(net),
    .B(n_3636_o_0),
    .C(n_3682_o_0),
    .Y(n_3683_o_0));
 AOI21xp33_ASAP7_75t_R n_3684 (.A1(n_3659_o_0),
    .A2(net86),
    .B(n_3683_o_0),
    .Y(n_3684_o_0));
 INVx1_ASAP7_75t_R n_3685 (.A(n_3673_o_0),
    .Y(n_3685_o_0));
 NAND2xp5_ASAP7_75t_R n_3686 (.A(n_3683_o_0),
    .B(n_3685_o_0),
    .Y(n_3686_o_0));
 INVx1_ASAP7_75t_R n_3687 (.A(n_3686_o_0),
    .Y(n_3687_o_0));
 OAI22xp33_ASAP7_75t_R n_3688 (.A1(n_3662_o_0),
    .A2(n_3680_o_0),
    .B1(n_3684_o_0),
    .B2(n_3687_o_0),
    .Y(n_3688_o_0));
 NOR3xp33_ASAP7_75t_R n_3689 (.A(n_3662_o_0),
    .B(n_3624_o_0),
    .C(n_3680_o_0),
    .Y(n_3689_o_0));
 XNOR2xp5_ASAP7_75t_R n_3690 (.A(_01047_),
    .B(_01051_),
    .Y(n_3690_o_0));
 XNOR2xp5_ASAP7_75t_R n_3691 (.A(_01087_),
    .B(_01095_),
    .Y(n_3691_o_0));
 XOR2xp5_ASAP7_75t_R n_3692 (.A(n_3690_o_0),
    .B(n_3691_o_0),
    .Y(n_3692_o_0));
 XNOR2xp5_ASAP7_75t_R n_3693 (.A(_01007_),
    .B(_01011_),
    .Y(n_3693_o_0));
 NAND2xp33_ASAP7_75t_R n_3694 (.A(_01048_),
    .B(n_3693_o_0),
    .Y(n_3694_o_0));
 OAI21xp33_ASAP7_75t_R n_3695 (.A1(_01048_),
    .A2(n_3693_o_0),
    .B(n_3694_o_0),
    .Y(n_3695_o_0));
 OAI21xp33_ASAP7_75t_R n_3696 (.A1(n_3695_o_0),
    .A2(n_3692_o_0),
    .B(net39),
    .Y(n_3696_o_0));
 AOI21xp33_ASAP7_75t_R n_3697 (.A1(n_3692_o_0),
    .A2(n_3695_o_0),
    .B(n_3696_o_0),
    .Y(n_3697_o_0));
 AOI21xp33_ASAP7_75t_R n_3698 (.A1(net3),
    .A2(_00672_),
    .B(n_3697_o_0),
    .Y(n_3698_o_0));
 NAND2xp33_ASAP7_75t_R n_3699 (.A(_00920_),
    .B(n_3698_o_0),
    .Y(n_3699_o_0));
 OAI21xp5_ASAP7_75t_R n_3700 (.A1(_00920_),
    .A2(n_3698_o_0),
    .B(n_3699_o_0),
    .Y(n_3700_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3701 (.A1(n_3624_o_0),
    .A2(n_3688_o_0),
    .B(n_3689_o_0),
    .C(n_3700_o_0),
    .Y(n_3701_o_0));
 XOR2xp5_ASAP7_75t_R n_3702 (.A(_00920_),
    .B(n_3698_o_0),
    .Y(n_3702_o_0));
 AO21x1_ASAP7_75t_R n_3703 (.A1(n_3635_o_0),
    .A2(n_3633_o_0),
    .B(n_2463_o_0),
    .Y(n_3703_o_0));
 OAI21xp33_ASAP7_75t_R n_3704 (.A1(net2),
    .A2(n_3638_o_0),
    .B(n_3674_o_0),
    .Y(n_3704_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3705 (.A1(net2),
    .A2(_00502_),
    .B(n_3703_o_0),
    .C(n_3704_o_0),
    .Y(n_3705_o_0));
 AOI21xp33_ASAP7_75t_R n_3706 (.A1(n_3645_o_0),
    .A2(n_3648_o_0),
    .B(n_3656_o_0),
    .Y(n_3706_o_0));
 AOI21xp33_ASAP7_75t_R n_3707 (.A1(net),
    .A2(n_3706_o_0),
    .B(n_3651_o_0),
    .Y(n_3707_o_0));
 NOR3xp33_ASAP7_75t_R n_3708 (.A(n_3705_o_0),
    .B(n_3707_o_0),
    .C(n_3658_o_0),
    .Y(n_3708_o_0));
 INVx1_ASAP7_75t_R n_3709 (.A(n_3637_o_0),
    .Y(n_3709_o_0));
 OAI22xp33_ASAP7_75t_R n_3710 (.A1(n_3709_o_0),
    .A2(n_3682_o_0),
    .B1(net25),
    .B2(net74),
    .Y(n_3710_o_0));
 INVx1_ASAP7_75t_R n_3711 (.A(n_3710_o_0),
    .Y(n_3711_o_0));
 NAND3xp33_ASAP7_75t_R n_3712 (.A(n_3642_o_0),
    .B(n_3659_o_0),
    .C(net50),
    .Y(n_3712_o_0));
 NAND3xp33_ASAP7_75t_R n_3713 (.A(n_3712_o_0),
    .B(n_3686_o_0),
    .C(n_3624_o_0),
    .Y(n_3713_o_0));
 OAI31xp33_ASAP7_75t_R n_3714 (.A1(n_3708_o_0),
    .A2(net41),
    .A3(n_3711_o_0),
    .B(n_3713_o_0),
    .Y(n_3714_o_0));
 XOR2xp5_ASAP7_75t_R n_3715 (.A(_01009_),
    .B(_01049_),
    .Y(n_3715_o_0));
 XNOR2xp5_ASAP7_75t_R n_3716 (.A(_01050_),
    .B(_01089_),
    .Y(n_3716_o_0));
 XNOR2xp5_ASAP7_75t_R n_3717 (.A(_01097_),
    .B(n_3716_o_0),
    .Y(n_3717_o_0));
 NOR2xp33_ASAP7_75t_R n_3718 (.A(n_3715_o_0),
    .B(n_3717_o_0),
    .Y(n_3718_o_0));
 NOR2xp33_ASAP7_75t_R n_3719 (.A(_00670_),
    .B(net),
    .Y(n_3719_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3720 (.A1(n_3715_o_0),
    .A2(n_3717_o_0),
    .B(n_3718_o_0),
    .C(net),
    .D(n_3719_o_0),
    .Y(n_3720_o_0));
 NOR2xp33_ASAP7_75t_R n_3721 (.A(_00922_),
    .B(n_3720_o_0),
    .Y(n_3721_o_0));
 AND2x2_ASAP7_75t_R n_3722 (.A(_00922_),
    .B(n_3720_o_0),
    .Y(n_3722_o_0));
 NOR2xp33_ASAP7_75t_R n_3723 (.A(n_3721_o_0),
    .B(n_3722_o_0),
    .Y(n_3723_o_0));
 INVx1_ASAP7_75t_R n_3724 (.A(n_3723_o_0),
    .Y(n_3724_o_0));
 AOI21xp33_ASAP7_75t_R n_3725 (.A1(n_3702_o_0),
    .A2(n_3714_o_0),
    .B(n_3724_o_0),
    .Y(n_3725_o_0));
 NOR2xp33_ASAP7_75t_R n_3726 (.A(_00500_),
    .B(net),
    .Y(n_3726_o_0));
 AOI21xp33_ASAP7_75t_R n_3727 (.A1(n_3666_o_0),
    .A2(n_3665_o_0),
    .B(n_3668_o_0),
    .Y(n_3727_o_0));
 INVx1_ASAP7_75t_R n_3728 (.A(n_3669_o_0),
    .Y(n_3728_o_0));
 OAI21xp33_ASAP7_75t_R n_3729 (.A1(n_3727_o_0),
    .A2(n_3728_o_0),
    .B(net),
    .Y(n_3729_o_0));
 INVx1_ASAP7_75t_R n_3730 (.A(n_3729_o_0),
    .Y(n_3730_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3731 (.A1(n_3670_o_0),
    .A2(net),
    .B(n_3671_o_0),
    .C(n_2421_o_0),
    .Y(n_3731_o_0));
 OAI311xp33_ASAP7_75t_R n_3732 (.A1(n_3726_o_0),
    .A2(n_3730_o_0),
    .A3(n_2421_o_0),
    .B1(n_3731_o_0),
    .C1(n_3659_o_0),
    .Y(n_3732_o_0));
 INVx1_ASAP7_75t_R n_3733 (.A(n_3726_o_0),
    .Y(n_3733_o_0));
 AOI21xp33_ASAP7_75t_R n_3734 (.A1(n_3733_o_0),
    .A2(n_3729_o_0),
    .B(_00916_),
    .Y(n_3734_o_0));
 OAI22xp33_ASAP7_75t_R n_3735 (.A1(n_3707_o_0),
    .A2(n_3658_o_0),
    .B1(n_3672_o_0),
    .B2(n_3734_o_0),
    .Y(n_3735_o_0));
 AOI22xp33_ASAP7_75t_R n_3736 (.A1(n_3732_o_0),
    .A2(n_3735_o_0),
    .B1(n_3641_o_0),
    .B2(n_3637_o_0),
    .Y(n_3736_o_0));
 NOR3xp33_ASAP7_75t_R n_3737 (.A(n_3705_o_0),
    .B(net74),
    .C(net50),
    .Y(n_3737_o_0));
 NOR2xp33_ASAP7_75t_R n_3738 (.A(n_3659_o_0),
    .B(n_3673_o_0),
    .Y(n_3738_o_0));
 INVx1_ASAP7_75t_R n_3739 (.A(n_3738_o_0),
    .Y(n_3739_o_0));
 AO21x1_ASAP7_75t_R n_3740 (.A1(n_3620_o_0),
    .A2(net),
    .B(n_3621_o_0),
    .Y(n_3740_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3741 (.A1(n_3620_o_0),
    .A2(net),
    .B(n_3621_o_0),
    .C(n_2399_o_0),
    .Y(n_3741_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3742 (.A1(n_2399_o_0),
    .A2(n_3740_o_0),
    .B(n_3741_o_0),
    .C(n_3683_o_0),
    .Y(n_3742_o_0));
 NAND2xp33_ASAP7_75t_R n_3743 (.A(n_3637_o_0),
    .B(n_3641_o_0),
    .Y(n_3743_o_0));
 AOI21xp33_ASAP7_75t_R n_3744 (.A1(net86),
    .A2(n_3660_o_0),
    .B(n_3743_o_0),
    .Y(n_3744_o_0));
 AOI22xp33_ASAP7_75t_R n_3745 (.A1(n_3739_o_0),
    .A2(n_3742_o_0),
    .B1(n_3627_o_0),
    .B2(n_3744_o_0),
    .Y(n_3745_o_0));
 OAI31xp33_ASAP7_75t_R n_3746 (.A1(net94),
    .A2(n_3736_o_0),
    .A3(n_3737_o_0),
    .B(n_3745_o_0),
    .Y(n_3746_o_0));
 XNOR2xp5_ASAP7_75t_R n_3747 (.A(_00922_),
    .B(n_3720_o_0),
    .Y(n_3747_o_0));
 INVx1_ASAP7_75t_R n_3748 (.A(n_3747_o_0),
    .Y(n_3748_o_0));
 AOI21xp33_ASAP7_75t_R n_3749 (.A1(n_3702_o_0),
    .A2(n_3746_o_0),
    .B(n_3748_o_0),
    .Y(n_3749_o_0));
 OAI211xp5_ASAP7_75t_R n_3750 (.A1(n_3682_o_0),
    .A2(n_3709_o_0),
    .B(n_3732_o_0),
    .C(n_3735_o_0),
    .Y(n_3750_o_0));
 NAND2xp33_ASAP7_75t_R n_3751 (.A(n_3627_o_0),
    .B(n_3750_o_0),
    .Y(n_3751_o_0));
 OAI211xp5_ASAP7_75t_R n_3752 (.A1(_00500_),
    .A2(net),
    .B(n_3729_o_0),
    .C(_00916_),
    .Y(n_3752_o_0));
 AOI22xp33_ASAP7_75t_R n_3753 (.A1(n_3752_o_0),
    .A2(n_3731_o_0),
    .B1(n_3678_o_0),
    .B2(n_3677_o_0),
    .Y(n_3753_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_3754 (.A1(net25),
    .A2(net74),
    .B(n_3753_o_0),
    .C(n_3676_o_0),
    .D(n_3623_o_0),
    .Y(n_3754_o_0));
 INVx1_ASAP7_75t_R n_3755 (.A(n_3754_o_0),
    .Y(n_3755_o_0));
 XNOR2xp5_ASAP7_75t_R n_3756 (.A(_00920_),
    .B(n_3698_o_0),
    .Y(n_3756_o_0));
 OAI211xp5_ASAP7_75t_R n_3757 (.A1(n_3751_o_0),
    .A2(n_3708_o_0),
    .B(n_3755_o_0),
    .C(n_3756_o_0),
    .Y(n_3757_o_0));
 AOI22xp33_ASAP7_75t_R n_3758 (.A1(n_3701_o_0),
    .A2(n_3725_o_0),
    .B1(n_3749_o_0),
    .B2(n_3757_o_0),
    .Y(n_3758_o_0));
 AOI21xp33_ASAP7_75t_R n_3759 (.A1(n_3623_o_0),
    .A2(n_3737_o_0),
    .B(n_3756_o_0),
    .Y(n_3759_o_0));
 INVx1_ASAP7_75t_R n_3760 (.A(n_3759_o_0),
    .Y(n_3760_o_0));
 NAND3xp33_ASAP7_75t_R n_3761 (.A(n_3685_o_0),
    .B(n_3642_o_0),
    .C(net74),
    .Y(n_3761_o_0));
 OAI21xp33_ASAP7_75t_R n_3762 (.A1(net50),
    .A2(n_3660_o_0),
    .B(n_3676_o_0),
    .Y(n_3762_o_0));
 NAND3xp33_ASAP7_75t_R n_3763 (.A(n_3761_o_0),
    .B(n_3762_o_0),
    .C(n_3627_o_0),
    .Y(n_3763_o_0));
 INVx1_ASAP7_75t_R n_3764 (.A(n_3763_o_0),
    .Y(n_3764_o_0));
 OAI21xp33_ASAP7_75t_R n_3765 (.A1(net86),
    .A2(n_3659_o_0),
    .B(n_3642_o_0),
    .Y(n_3765_o_0));
 NAND2xp33_ASAP7_75t_R n_3766 (.A(net50),
    .B(n_3683_o_0),
    .Y(n_3766_o_0));
 AOI21xp33_ASAP7_75t_R n_3767 (.A1(n_3765_o_0),
    .A2(n_3766_o_0),
    .B(n_3627_o_0),
    .Y(n_3767_o_0));
 NAND2xp33_ASAP7_75t_R n_3768 (.A(net30),
    .B(n_3642_o_0),
    .Y(n_3768_o_0));
 AOI211xp5_ASAP7_75t_R n_3769 (.A1(net50),
    .A2(n_3659_o_0),
    .B(n_3753_o_0),
    .C(n_3705_o_0),
    .Y(n_3769_o_0));
 INVx1_ASAP7_75t_R n_3770 (.A(n_3700_o_0),
    .Y(n_3770_o_0));
 AOI21xp33_ASAP7_75t_R n_3771 (.A1(net93),
    .A2(n_3769_o_0),
    .B(n_3770_o_0),
    .Y(n_3771_o_0));
 OAI21xp33_ASAP7_75t_R n_3772 (.A1(n_3627_o_0),
    .A2(n_3768_o_0),
    .B(n_3771_o_0),
    .Y(n_3772_o_0));
 OAI31xp33_ASAP7_75t_R n_3773 (.A1(n_3760_o_0),
    .A2(n_3764_o_0),
    .A3(n_3767_o_0),
    .B(n_3772_o_0),
    .Y(n_3773_o_0));
 NOR3xp33_ASAP7_75t_R n_3774 (.A(n_3685_o_0),
    .B(net72),
    .C(net30),
    .Y(n_3774_o_0));
 NOR4xp25_ASAP7_75t_R n_3775 (.A(n_3707_o_0),
    .B(n_3658_o_0),
    .C(n_3672_o_0),
    .D(n_3734_o_0),
    .Y(n_3775_o_0));
 OAI22xp33_ASAP7_75t_R n_3776 (.A1(n_3775_o_0),
    .A2(n_3753_o_0),
    .B1(n_3682_o_0),
    .B2(n_3709_o_0),
    .Y(n_3776_o_0));
 AO22x1_ASAP7_75t_R n_3777 (.A1(n_3627_o_0),
    .A2(n_3774_o_0),
    .B1(n_3776_o_0),
    .B2(n_3624_o_0),
    .Y(n_3777_o_0));
 NOR2xp33_ASAP7_75t_R n_3778 (.A(n_3673_o_0),
    .B(n_3660_o_0),
    .Y(n_3778_o_0));
 INVx1_ASAP7_75t_R n_3779 (.A(n_3778_o_0),
    .Y(n_3779_o_0));
 NAND4xp25_ASAP7_75t_R n_3780 (.A(n_3712_o_0),
    .B(n_3686_o_0),
    .C(n_3702_o_0),
    .D(n_3624_o_0),
    .Y(n_3780_o_0));
 OAI311xp33_ASAP7_75t_R n_3781 (.A1(n_3624_o_0),
    .A2(n_3705_o_0),
    .A3(n_3779_o_0),
    .B1(n_3723_o_0),
    .C1(n_3780_o_0),
    .Y(n_3781_o_0));
 INVx1_ASAP7_75t_R n_3782 (.A(n_3613_o_0),
    .Y(n_3782_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3783 (.A1(n_3700_o_0),
    .A2(n_3777_o_0),
    .B(n_3781_o_0),
    .C(n_3782_o_0),
    .Y(n_3783_o_0));
 AOI21xp33_ASAP7_75t_R n_3784 (.A1(n_3747_o_0),
    .A2(n_3773_o_0),
    .B(n_3783_o_0),
    .Y(n_3784_o_0));
 AOI21xp33_ASAP7_75t_R n_3785 (.A1(n_3613_o_0),
    .A2(n_3758_o_0),
    .B(n_3784_o_0),
    .Y(n_3785_o_0));
 NOR2xp33_ASAP7_75t_R n_3786 (.A(n_3673_o_0),
    .B(n_3683_o_0),
    .Y(n_3786_o_0));
 INVx1_ASAP7_75t_R n_3787 (.A(n_3786_o_0),
    .Y(n_3787_o_0));
 AOI21xp33_ASAP7_75t_R n_3788 (.A1(n_3685_o_0),
    .A2(n_3708_o_0),
    .B(net90),
    .Y(n_3788_o_0));
 NAND2xp33_ASAP7_75t_R n_3789 (.A(n_3659_o_0),
    .B(n_3673_o_0),
    .Y(n_3789_o_0));
 INVx1_ASAP7_75t_R n_3790 (.A(n_3789_o_0),
    .Y(n_3790_o_0));
 OAI21xp33_ASAP7_75t_R n_3791 (.A1(n_3743_o_0),
    .A2(n_3790_o_0),
    .B(net90),
    .Y(n_3791_o_0));
 OAI21xp33_ASAP7_75t_R n_3792 (.A1(n_3736_o_0),
    .A2(n_3791_o_0),
    .B(n_3756_o_0),
    .Y(n_3792_o_0));
 AOI21xp33_ASAP7_75t_R n_3793 (.A1(n_3787_o_0),
    .A2(n_3788_o_0),
    .B(n_3792_o_0),
    .Y(n_3793_o_0));
 AOI22xp33_ASAP7_75t_R n_3794 (.A1(n_3685_o_0),
    .A2(n_3659_o_0),
    .B1(n_3637_o_0),
    .B2(n_3641_o_0),
    .Y(n_3794_o_0));
 OAI31xp33_ASAP7_75t_R n_3795 (.A1(net11),
    .A2(n_3680_o_0),
    .A3(n_3794_o_0),
    .B(n_3770_o_0),
    .Y(n_3795_o_0));
 AOI21xp33_ASAP7_75t_R n_3796 (.A1(n_3686_o_0),
    .A2(n_3627_o_0),
    .B(n_3795_o_0),
    .Y(n_3796_o_0));
 OAI31xp33_ASAP7_75t_R n_3797 (.A1(n_3747_o_0),
    .A2(n_3793_o_0),
    .A3(n_3796_o_0),
    .B(n_3613_o_0),
    .Y(n_3797_o_0));
 NOR2xp33_ASAP7_75t_R n_3798 (.A(n_3659_o_0),
    .B(n_3673_o_0),
    .Y(n_3798_o_0));
 INVx1_ASAP7_75t_R n_3799 (.A(n_3798_o_0),
    .Y(n_3799_o_0));
 AOI21xp33_ASAP7_75t_R n_3800 (.A1(n_3642_o_0),
    .A2(net86),
    .B(n_3626_o_0),
    .Y(n_3800_o_0));
 NAND2xp33_ASAP7_75t_R n_3801 (.A(net50),
    .B(n_3642_o_0),
    .Y(n_3801_o_0));
 AOI21xp33_ASAP7_75t_R n_3802 (.A1(n_3801_o_0),
    .A2(n_3799_o_0),
    .B(n_3627_o_0),
    .Y(n_3802_o_0));
 AOI21xp33_ASAP7_75t_R n_3803 (.A1(n_3799_o_0),
    .A2(n_3800_o_0),
    .B(n_3802_o_0),
    .Y(n_3803_o_0));
 NOR2xp33_ASAP7_75t_R n_3804 (.A(n_3626_o_0),
    .B(n_3736_o_0),
    .Y(n_3804_o_0));
 NAND4xp25_ASAP7_75t_R n_3805 (.A(n_3676_o_0),
    .B(net50),
    .C(n_3678_o_0),
    .D(n_3677_o_0),
    .Y(n_3805_o_0));
 OAI21xp33_ASAP7_75t_R n_3806 (.A1(net74),
    .A2(n_3685_o_0),
    .B(n_3642_o_0),
    .Y(n_3806_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3807 (.A1(n_3642_o_0),
    .A2(n_3738_o_0),
    .B(n_3806_o_0),
    .C(n_3627_o_0),
    .Y(n_3807_o_0));
 AOI211xp5_ASAP7_75t_R n_3808 (.A1(n_3804_o_0),
    .A2(n_3805_o_0),
    .B(n_3756_o_0),
    .C(n_3807_o_0),
    .Y(n_3808_o_0));
 AOI211xp5_ASAP7_75t_R n_3809 (.A1(n_3700_o_0),
    .A2(n_3803_o_0),
    .B(n_3808_o_0),
    .C(n_3748_o_0),
    .Y(n_3809_o_0));
 INVx1_ASAP7_75t_R n_3810 (.A(n_3742_o_0),
    .Y(n_3810_o_0));
 OAI211xp5_ASAP7_75t_R n_3811 (.A1(n_3685_o_0),
    .A2(net74),
    .B(n_3637_o_0),
    .C(n_3641_o_0),
    .Y(n_3811_o_0));
 AOI31xp33_ASAP7_75t_R n_3812 (.A1(net90),
    .A2(n_3811_o_0),
    .A3(n_3761_o_0),
    .B(n_3700_o_0),
    .Y(n_3812_o_0));
 OAI21xp33_ASAP7_75t_R n_3813 (.A1(n_3739_o_0),
    .A2(n_3810_o_0),
    .B(n_3812_o_0),
    .Y(n_3813_o_0));
 NAND2xp33_ASAP7_75t_R n_3814 (.A(n_3642_o_0),
    .B(n_3738_o_0),
    .Y(n_3814_o_0));
 NAND3xp33_ASAP7_75t_R n_3815 (.A(n_3660_o_0),
    .B(n_3676_o_0),
    .C(net86),
    .Y(n_3815_o_0));
 AOI31xp33_ASAP7_75t_R n_3816 (.A1(n_3627_o_0),
    .A2(n_3761_o_0),
    .A3(n_3815_o_0),
    .B(n_3702_o_0),
    .Y(n_3816_o_0));
 OAI21xp33_ASAP7_75t_R n_3817 (.A1(n_3814_o_0),
    .A2(net94),
    .B(n_3816_o_0),
    .Y(n_3817_o_0));
 NAND3xp33_ASAP7_75t_R n_3818 (.A(n_3813_o_0),
    .B(n_3817_o_0),
    .C(n_3724_o_0),
    .Y(n_3818_o_0));
 OAI21xp33_ASAP7_75t_R n_3819 (.A1(n_3811_o_0),
    .A2(net94),
    .B(n_3770_o_0),
    .Y(n_3819_o_0));
 OAI21xp33_ASAP7_75t_R n_3820 (.A1(net50),
    .A2(n_3659_o_0),
    .B(n_3732_o_0),
    .Y(n_3820_o_0));
 AOI21xp33_ASAP7_75t_R n_3821 (.A1(n_3642_o_0),
    .A2(net74),
    .B(n_3626_o_0),
    .Y(n_3821_o_0));
 OAI21xp33_ASAP7_75t_R n_3822 (.A1(n_3705_o_0),
    .A2(n_3820_o_0),
    .B(n_3821_o_0),
    .Y(n_3822_o_0));
 OAI31xp33_ASAP7_75t_R n_3823 (.A1(net94),
    .A2(net72),
    .A3(n_3685_o_0),
    .B(n_3822_o_0),
    .Y(n_3823_o_0));
 OAI21xp33_ASAP7_75t_R n_3824 (.A1(n_3705_o_0),
    .A2(n_3739_o_0),
    .B(n_3627_o_0),
    .Y(n_3824_o_0));
 OA21x2_ASAP7_75t_R n_3825 (.A1(n_3794_o_0),
    .A2(net63),
    .B(n_3756_o_0),
    .Y(n_3825_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3826 (.A1(n_3824_o_0),
    .A2(n_3711_o_0),
    .B(n_3825_o_0),
    .C(n_3747_o_0),
    .Y(n_3826_o_0));
 OAI21xp33_ASAP7_75t_R n_3827 (.A1(n_3819_o_0),
    .A2(n_3823_o_0),
    .B(n_3826_o_0),
    .Y(n_3827_o_0));
 XNOR2xp5_ASAP7_75t_R n_3828 (.A(_00921_),
    .B(n_3602_o_0),
    .Y(n_3828_o_0));
 AOI31xp33_ASAP7_75t_R n_3829 (.A1(n_3782_o_0),
    .A2(n_3818_o_0),
    .A3(n_3827_o_0),
    .B(n_3828_o_0),
    .Y(n_3829_o_0));
 OAI21xp33_ASAP7_75t_R n_3830 (.A1(n_3797_o_0),
    .A2(n_3809_o_0),
    .B(n_3829_o_0),
    .Y(n_3830_o_0));
 OAI21xp33_ASAP7_75t_R n_3831 (.A1(n_3605_o_0),
    .A2(n_3785_o_0),
    .B(n_3830_o_0),
    .Y(n_3831_o_0));
 NOR2xp33_ASAP7_75t_R n_3832 (.A(n_3623_o_0),
    .B(n_3736_o_0),
    .Y(n_3832_o_0));
 INVx1_ASAP7_75t_R n_3833 (.A(n_3832_o_0),
    .Y(n_3833_o_0));
 AOI31xp33_ASAP7_75t_R n_3834 (.A1(n_3686_o_0),
    .A2(n_3712_o_0),
    .A3(n_3627_o_0),
    .B(n_3700_o_0),
    .Y(n_3834_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3835 (.A1(net25),
    .A2(net30),
    .B(net72),
    .C(n_3627_o_0),
    .Y(n_3835_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3836 (.A1(n_3676_o_0),
    .A2(n_3739_o_0),
    .B(n_3835_o_0),
    .C(n_3756_o_0),
    .Y(n_3836_o_0));
 AOI31xp33_ASAP7_75t_R n_3837 (.A1(n_3624_o_0),
    .A2(n_3750_o_0),
    .A3(n_3805_o_0),
    .B(n_3836_o_0),
    .Y(n_3837_o_0));
 AOI211xp5_ASAP7_75t_R n_3838 (.A1(n_3833_o_0),
    .A2(n_3834_o_0),
    .B(n_3837_o_0),
    .C(n_3605_o_0),
    .Y(n_3838_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3839 (.A1(n_3739_o_0),
    .A2(n_3642_o_0),
    .B(n_3769_o_0),
    .C(net41),
    .Y(n_3839_o_0));
 AOI31xp33_ASAP7_75t_R n_3840 (.A1(net25),
    .A2(net72),
    .A3(n_3627_o_0),
    .B(n_3702_o_0),
    .Y(n_3840_o_0));
 OA21x2_ASAP7_75t_R n_3841 (.A1(n_3739_o_0),
    .A2(n_3810_o_0),
    .B(n_3840_o_0),
    .Y(n_3841_o_0));
 INVx1_ASAP7_75t_R n_3842 (.A(n_3737_o_0),
    .Y(n_3842_o_0));
 AOI21xp33_ASAP7_75t_R n_3843 (.A1(n_3660_o_0),
    .A2(n_3683_o_0),
    .B(n_3623_o_0),
    .Y(n_3843_o_0));
 INVx1_ASAP7_75t_R n_3844 (.A(n_3843_o_0),
    .Y(n_3844_o_0));
 OAI21xp33_ASAP7_75t_R n_3845 (.A1(n_3794_o_0),
    .A2(n_3844_o_0),
    .B(n_3770_o_0),
    .Y(n_3845_o_0));
 INVx1_ASAP7_75t_R n_3846 (.A(n_3828_o_0),
    .Y(n_3846_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3847 (.A1(n_3842_o_0),
    .A2(n_3800_o_0),
    .B(n_3845_o_0),
    .C(n_3846_o_0),
    .Y(n_3847_o_0));
 AOI21xp33_ASAP7_75t_R n_3848 (.A1(n_3839_o_0),
    .A2(n_3841_o_0),
    .B(n_3847_o_0),
    .Y(n_3848_o_0));
 NOR3xp33_ASAP7_75t_R n_3849 (.A(n_3838_o_0),
    .B(n_3848_o_0),
    .C(n_3724_o_0),
    .Y(n_3849_o_0));
 NOR2xp33_ASAP7_75t_R n_3850 (.A(net30),
    .B(n_3642_o_0),
    .Y(n_3850_o_0));
 NAND3xp33_ASAP7_75t_R n_3851 (.A(n_3815_o_0),
    .B(n_3712_o_0),
    .C(n_3627_o_0),
    .Y(n_3851_o_0));
 OAI31xp33_ASAP7_75t_R n_3852 (.A1(n_3605_o_0),
    .A2(net94),
    .A3(n_3850_o_0),
    .B(n_3851_o_0),
    .Y(n_3852_o_0));
 OAI21xp33_ASAP7_75t_R n_3853 (.A1(n_3794_o_0),
    .A2(n_3844_o_0),
    .B(n_3828_o_0),
    .Y(n_3853_o_0));
 AOI21xp33_ASAP7_75t_R n_3854 (.A1(n_3679_o_0),
    .A2(n_3800_o_0),
    .B(n_3853_o_0),
    .Y(n_3854_o_0));
 NAND2xp33_ASAP7_75t_R n_3855 (.A(net74),
    .B(net50),
    .Y(n_3855_o_0));
 INVx1_ASAP7_75t_R n_3856 (.A(n_3855_o_0),
    .Y(n_3856_o_0));
 NOR3xp33_ASAP7_75t_R n_3857 (.A(n_3856_o_0),
    .B(net72),
    .C(net63),
    .Y(n_3857_o_0));
 NAND2xp33_ASAP7_75t_R n_3858 (.A(n_3659_o_0),
    .B(n_3685_o_0),
    .Y(n_3858_o_0));
 NOR2xp33_ASAP7_75t_R n_3859 (.A(n_3642_o_0),
    .B(n_3623_o_0),
    .Y(n_3859_o_0));
 AOI21xp33_ASAP7_75t_R n_3860 (.A1(n_3858_o_0),
    .A2(n_3859_o_0),
    .B(n_3604_o_0),
    .Y(n_3860_o_0));
 OAI21xp33_ASAP7_75t_R n_3861 (.A1(n_3786_o_0),
    .A2(n_3824_o_0),
    .B(n_3860_o_0),
    .Y(n_3861_o_0));
 OAI21xp33_ASAP7_75t_R n_3862 (.A1(n_3857_o_0),
    .A2(n_3861_o_0),
    .B(n_3700_o_0),
    .Y(n_3862_o_0));
 OAI21xp33_ASAP7_75t_R n_3863 (.A1(n_3854_o_0),
    .A2(n_3862_o_0),
    .B(n_3747_o_0),
    .Y(n_3863_o_0));
 AOI21xp33_ASAP7_75t_R n_3864 (.A1(n_3702_o_0),
    .A2(n_3852_o_0),
    .B(n_3863_o_0),
    .Y(n_3864_o_0));
 NAND3xp33_ASAP7_75t_R n_3865 (.A(n_3750_o_0),
    .B(n_3805_o_0),
    .C(n_3624_o_0),
    .Y(n_3865_o_0));
 OAI31xp33_ASAP7_75t_R n_3866 (.A1(net72),
    .A2(net41),
    .A3(n_3779_o_0),
    .B(n_3865_o_0),
    .Y(n_3866_o_0));
 OAI21xp33_ASAP7_75t_R n_3867 (.A1(n_3705_o_0),
    .A2(n_3820_o_0),
    .B(n_3627_o_0),
    .Y(n_3867_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3868 (.A1(n_3786_o_0),
    .A2(n_3856_o_0),
    .B(n_3624_o_0),
    .C(n_3846_o_0),
    .Y(n_3868_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3869 (.A1(n_3867_o_0),
    .A2(n_3786_o_0),
    .B(n_3868_o_0),
    .C(n_3747_o_0),
    .Y(n_3869_o_0));
 OA21x2_ASAP7_75t_R n_3870 (.A1(n_3604_o_0),
    .A2(n_3866_o_0),
    .B(n_3869_o_0),
    .Y(n_3870_o_0));
 OAI21xp33_ASAP7_75t_R n_3871 (.A1(n_3684_o_0),
    .A2(n_3755_o_0),
    .B(n_3828_o_0),
    .Y(n_3871_o_0));
 INVx1_ASAP7_75t_R n_3872 (.A(n_3821_o_0),
    .Y(n_3872_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3873 (.A1(n_3798_o_0),
    .A2(n_3872_o_0),
    .B(n_3860_o_0),
    .C(n_3723_o_0),
    .Y(n_3873_o_0));
 OA21x2_ASAP7_75t_R n_3874 (.A1(n_3764_o_0),
    .A2(n_3871_o_0),
    .B(n_3873_o_0),
    .Y(n_3874_o_0));
 NAND3xp33_ASAP7_75t_R n_3875 (.A(n_3778_o_0),
    .B(n_3676_o_0),
    .C(n_3623_o_0),
    .Y(n_3875_o_0));
 OAI21xp33_ASAP7_75t_R n_3876 (.A1(net63),
    .A2(n_3708_o_0),
    .B(n_3875_o_0),
    .Y(n_3876_o_0));
 AOI211xp5_ASAP7_75t_R n_3877 (.A1(n_3642_o_0),
    .A2(n_3660_o_0),
    .B(n_3876_o_0),
    .C(n_3846_o_0),
    .Y(n_3877_o_0));
 INVx1_ASAP7_75t_R n_3878 (.A(n_3766_o_0),
    .Y(n_3878_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3879 (.A1(n_3641_o_0),
    .A2(n_3637_o_0),
    .B(n_3778_o_0),
    .C(n_3627_o_0),
    .Y(n_3879_o_0));
 OAI21xp33_ASAP7_75t_R n_3880 (.A1(n_3878_o_0),
    .A2(n_3879_o_0),
    .B(n_3605_o_0),
    .Y(n_3880_o_0));
 AOI21xp33_ASAP7_75t_R n_3881 (.A1(n_3832_o_0),
    .A2(n_3686_o_0),
    .B(n_3880_o_0),
    .Y(n_3881_o_0));
 NAND2xp33_ASAP7_75t_R n_3882 (.A(n_3683_o_0),
    .B(n_3789_o_0),
    .Y(n_3882_o_0));
 OAI311xp33_ASAP7_75t_R n_3883 (.A1(net72),
    .A2(net30),
    .A3(n_3742_o_0),
    .B1(n_3624_o_0),
    .C1(n_3882_o_0),
    .Y(n_3883_o_0));
 NAND3xp33_ASAP7_75t_R n_3884 (.A(n_3742_o_0),
    .B(n_3855_o_0),
    .C(net63),
    .Y(n_3884_o_0));
 AOI211xp5_ASAP7_75t_R n_3885 (.A1(n_3883_o_0),
    .A2(n_3884_o_0),
    .B(n_3604_o_0),
    .C(n_3747_o_0),
    .Y(n_3885_o_0));
 NOR2xp33_ASAP7_75t_R n_3886 (.A(n_3747_o_0),
    .B(n_3605_o_0),
    .Y(n_3886_o_0));
 AOI211xp5_ASAP7_75t_R n_3887 (.A1(n_3778_o_0),
    .A2(n_3676_o_0),
    .B(net93),
    .C(n_3736_o_0),
    .Y(n_3887_o_0));
 AOI31xp33_ASAP7_75t_R n_3888 (.A1(n_3627_o_0),
    .A2(n_3765_o_0),
    .A3(n_3766_o_0),
    .B(n_3887_o_0),
    .Y(n_3888_o_0));
 OAI22xp33_ASAP7_75t_R n_3889 (.A1(n_3885_o_0),
    .A2(n_3886_o_0),
    .B1(n_3888_o_0),
    .B2(n_3605_o_0),
    .Y(n_3889_o_0));
 OAI31xp33_ASAP7_75t_R n_3890 (.A1(n_3723_o_0),
    .A2(n_3877_o_0),
    .A3(n_3881_o_0),
    .B(n_3889_o_0),
    .Y(n_3890_o_0));
 OAI321xp33_ASAP7_75t_R n_3891 (.A1(n_3700_o_0),
    .A2(n_3870_o_0),
    .A3(n_3874_o_0),
    .B1(n_3890_o_0),
    .B2(n_3702_o_0),
    .C(n_3782_o_0),
    .Y(n_3891_o_0));
 OAI31xp33_ASAP7_75t_R n_3892 (.A1(n_3782_o_0),
    .A2(n_3849_o_0),
    .A3(n_3864_o_0),
    .B(n_3891_o_0),
    .Y(n_3892_o_0));
 INVx1_ASAP7_75t_R n_3893 (.A(n_3882_o_0),
    .Y(n_3893_o_0));
 NAND2xp33_ASAP7_75t_R n_3894 (.A(net74),
    .B(n_3642_o_0),
    .Y(n_3894_o_0));
 OAI211xp5_ASAP7_75t_R n_3895 (.A1(n_3679_o_0),
    .A2(net25),
    .B(n_3894_o_0),
    .C(n_3624_o_0),
    .Y(n_3895_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3896 (.A1(n_3893_o_0),
    .A2(n_3879_o_0),
    .B(n_3895_o_0),
    .C(n_3770_o_0),
    .Y(n_3896_o_0));
 INVx1_ASAP7_75t_R n_3897 (.A(n_3822_o_0),
    .Y(n_3897_o_0));
 AOI21xp33_ASAP7_75t_R n_3898 (.A1(n_3762_o_0),
    .A2(n_3761_o_0),
    .B(n_3627_o_0),
    .Y(n_3898_o_0));
 OAI31xp33_ASAP7_75t_R n_3899 (.A1(n_3756_o_0),
    .A2(n_3897_o_0),
    .A3(n_3898_o_0),
    .B(n_3604_o_0),
    .Y(n_3899_o_0));
 INVx1_ASAP7_75t_R n_3900 (.A(n_3801_o_0),
    .Y(n_3900_o_0));
 OAI311xp33_ASAP7_75t_R n_3901 (.A1(n_3682_o_0),
    .A2(n_3709_o_0),
    .A3(net30),
    .B1(n_3627_o_0),
    .C1(n_3750_o_0),
    .Y(n_3901_o_0));
 OAI31xp33_ASAP7_75t_R n_3902 (.A1(net11),
    .A2(n_3900_o_0),
    .A3(n_3737_o_0),
    .B(n_3901_o_0),
    .Y(n_3902_o_0));
 AOI21xp33_ASAP7_75t_R n_3903 (.A1(net25),
    .A2(n_3708_o_0),
    .B(n_3684_o_0),
    .Y(n_3903_o_0));
 AOI211xp5_ASAP7_75t_R n_3904 (.A1(n_3903_o_0),
    .A2(n_3624_o_0),
    .B(n_3700_o_0),
    .C(n_3788_o_0),
    .Y(n_3904_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3905 (.A1(n_3700_o_0),
    .A2(n_3902_o_0),
    .B(n_3904_o_0),
    .C(n_3605_o_0),
    .Y(n_3905_o_0));
 OAI21xp33_ASAP7_75t_R n_3906 (.A1(n_3896_o_0),
    .A2(n_3899_o_0),
    .B(n_3905_o_0),
    .Y(n_3906_o_0));
 NAND2xp33_ASAP7_75t_R n_3907 (.A(net30),
    .B(n_3624_o_0),
    .Y(n_3907_o_0));
 NAND2xp33_ASAP7_75t_R n_3908 (.A(n_3762_o_0),
    .B(n_3702_o_0),
    .Y(n_3908_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3909 (.A1(n_3642_o_0),
    .A2(n_3907_o_0),
    .B(n_3908_o_0),
    .C(n_3828_o_0),
    .Y(n_3909_o_0));
 NAND2xp33_ASAP7_75t_R n_3910 (.A(n_3676_o_0),
    .B(n_3778_o_0),
    .Y(n_3910_o_0));
 OAI21xp33_ASAP7_75t_R n_3911 (.A1(n_3642_o_0),
    .A2(n_3789_o_0),
    .B(n_3627_o_0),
    .Y(n_3911_o_0));
 AOI211xp5_ASAP7_75t_R n_3912 (.A1(n_3641_o_0),
    .A2(n_3637_o_0),
    .B(n_3685_o_0),
    .C(net74),
    .Y(n_3912_o_0));
 AOI22xp33_ASAP7_75t_R n_3913 (.A1(n_3911_o_0),
    .A2(n_3756_o_0),
    .B1(net63),
    .B2(n_3912_o_0),
    .Y(n_3913_o_0));
 AOI31xp33_ASAP7_75t_R n_3914 (.A1(n_3624_o_0),
    .A2(n_3801_o_0),
    .A3(n_3910_o_0),
    .B(n_3913_o_0),
    .Y(n_3914_o_0));
 AOI21xp33_ASAP7_75t_R n_3915 (.A1(n_3800_o_0),
    .A2(n_3815_o_0),
    .B(n_3700_o_0),
    .Y(n_3915_o_0));
 INVx1_ASAP7_75t_R n_3916 (.A(n_3915_o_0),
    .Y(n_3916_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3917 (.A1(n_3682_o_0),
    .A2(n_3709_o_0),
    .B(n_3685_o_0),
    .C(net30),
    .Y(n_3917_o_0));
 AOI31xp33_ASAP7_75t_R n_3918 (.A1(net25),
    .A2(n_3683_o_0),
    .A3(net30),
    .B(n_3626_o_0),
    .Y(n_3918_o_0));
 AOI21xp33_ASAP7_75t_R n_3919 (.A1(n_3801_o_0),
    .A2(n_3918_o_0),
    .B(n_3702_o_0),
    .Y(n_3919_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3920 (.A1(n_3917_o_0),
    .A2(net63),
    .B(n_3919_o_0),
    .C(n_3828_o_0),
    .Y(n_3920_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3921 (.A1(n_3750_o_0),
    .A2(n_3754_o_0),
    .B(n_3916_o_0),
    .C(n_3920_o_0),
    .Y(n_3921_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3922 (.A1(n_3909_o_0),
    .A2(n_3914_o_0),
    .B(n_3921_o_0),
    .C(n_3724_o_0),
    .Y(n_3922_o_0));
 AO21x1_ASAP7_75t_R n_3923 (.A1(n_3906_o_0),
    .A2(n_3747_o_0),
    .B(n_3922_o_0),
    .Y(n_3923_o_0));
 AOI211xp5_ASAP7_75t_R n_3924 (.A1(n_3642_o_0),
    .A2(net30),
    .B(n_3798_o_0),
    .C(net93),
    .Y(n_3924_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3925 (.A1(net30),
    .A2(n_3642_o_0),
    .B(n_3627_o_0),
    .C(n_3924_o_0),
    .Y(n_3925_o_0));
 INVx1_ASAP7_75t_R n_3926 (.A(n_3769_o_0),
    .Y(n_3926_o_0));
 AOI211xp5_ASAP7_75t_R n_3927 (.A1(net25),
    .A2(n_3683_o_0),
    .B(n_3626_o_0),
    .C(net30),
    .Y(n_3927_o_0));
 AOI31xp33_ASAP7_75t_R n_3928 (.A1(n_3624_o_0),
    .A2(n_3926_o_0),
    .A3(n_3806_o_0),
    .B(n_3927_o_0),
    .Y(n_3928_o_0));
 OAI21xp33_ASAP7_75t_R n_3929 (.A1(n_3770_o_0),
    .A2(n_3928_o_0),
    .B(n_3604_o_0),
    .Y(n_3929_o_0));
 OAI21xp33_ASAP7_75t_R n_3930 (.A1(n_3786_o_0),
    .A2(n_3844_o_0),
    .B(n_3756_o_0),
    .Y(n_3930_o_0));
 AOI21xp33_ASAP7_75t_R n_3931 (.A1(n_3761_o_0),
    .A2(n_3754_o_0),
    .B(n_3700_o_0),
    .Y(n_3931_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3932 (.A1(n_3768_o_0),
    .A2(net41),
    .B(n_3931_o_0),
    .C(n_3828_o_0),
    .Y(n_3932_o_0));
 OAI21xp33_ASAP7_75t_R n_3933 (.A1(n_3930_o_0),
    .A2(n_3897_o_0),
    .B(n_3932_o_0),
    .Y(n_3933_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3934 (.A1(n_3770_o_0),
    .A2(n_3925_o_0),
    .B(n_3929_o_0),
    .C(n_3933_o_0),
    .Y(n_3934_o_0));
 INVx1_ASAP7_75t_R n_3935 (.A(n_3762_o_0),
    .Y(n_3935_o_0));
 OAI31xp33_ASAP7_75t_R n_3936 (.A1(net11),
    .A2(n_3935_o_0),
    .A3(n_3736_o_0),
    .B(n_3770_o_0),
    .Y(n_3936_o_0));
 OAI21xp33_ASAP7_75t_R n_3937 (.A1(net25),
    .A2(net74),
    .B(n_3742_o_0),
    .Y(n_3937_o_0));
 INVx1_ASAP7_75t_R n_3938 (.A(n_3937_o_0),
    .Y(n_3938_o_0));
 INVx1_ASAP7_75t_R n_3939 (.A(n_3815_o_0),
    .Y(n_3939_o_0));
 INVx1_ASAP7_75t_R n_3940 (.A(n_3712_o_0),
    .Y(n_3940_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3941 (.A1(n_3682_o_0),
    .A2(n_3709_o_0),
    .B(net25),
    .C(n_3623_o_0),
    .Y(n_3941_o_0));
 AOI21xp33_ASAP7_75t_R n_3942 (.A1(n_3805_o_0),
    .A2(n_3941_o_0),
    .B(n_3702_o_0),
    .Y(n_3942_o_0));
 OAI31xp33_ASAP7_75t_R n_3943 (.A1(net41),
    .A2(n_3939_o_0),
    .A3(n_3940_o_0),
    .B(n_3942_o_0),
    .Y(n_3943_o_0));
 OAI211xp5_ASAP7_75t_R n_3944 (.A1(n_3936_o_0),
    .A2(n_3938_o_0),
    .B(n_3846_o_0),
    .C(n_3943_o_0),
    .Y(n_3944_o_0));
 OAI21xp33_ASAP7_75t_R n_3945 (.A1(net25),
    .A2(n_3679_o_0),
    .B(n_3627_o_0),
    .Y(n_3945_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3946 (.A1(n_3642_o_0),
    .A2(net30),
    .B(net11),
    .C(n_3945_o_0),
    .Y(n_3946_o_0));
 NAND3xp33_ASAP7_75t_R n_3947 (.A(net93),
    .B(net72),
    .C(net30),
    .Y(n_3947_o_0));
 AOI31xp33_ASAP7_75t_R n_3948 (.A1(n_3947_o_0),
    .A2(n_3895_o_0),
    .A3(n_3756_o_0),
    .B(n_3605_o_0),
    .Y(n_3948_o_0));
 OAI21xp33_ASAP7_75t_R n_3949 (.A1(n_3700_o_0),
    .A2(n_3946_o_0),
    .B(n_3948_o_0),
    .Y(n_3949_o_0));
 NAND3xp33_ASAP7_75t_R n_3950 (.A(n_3944_o_0),
    .B(n_3949_o_0),
    .C(n_3747_o_0),
    .Y(n_3950_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3951 (.A1(n_3724_o_0),
    .A2(n_3934_o_0),
    .B(n_3950_o_0),
    .C(n_3613_o_0),
    .Y(n_3951_o_0));
 AOI21xp33_ASAP7_75t_R n_3952 (.A1(n_3613_o_0),
    .A2(n_3923_o_0),
    .B(n_3951_o_0),
    .Y(n_3952_o_0));
 AOI211xp5_ASAP7_75t_R n_3953 (.A1(n_3804_o_0),
    .A2(n_3811_o_0),
    .B(n_3770_o_0),
    .C(n_3802_o_0),
    .Y(n_3953_o_0));
 INVx1_ASAP7_75t_R n_3954 (.A(n_3953_o_0),
    .Y(n_3954_o_0));
 NAND3xp33_ASAP7_75t_R n_3955 (.A(n_3843_o_0),
    .B(n_3806_o_0),
    .C(n_3766_o_0),
    .Y(n_3955_o_0));
 NAND4xp25_ASAP7_75t_R n_3956 (.A(n_3926_o_0),
    .B(n_3787_o_0),
    .C(n_3661_o_0),
    .D(n_3627_o_0),
    .Y(n_3956_o_0));
 AOI31xp33_ASAP7_75t_R n_3957 (.A1(n_3955_o_0),
    .A2(n_3956_o_0),
    .A3(n_3770_o_0),
    .B(n_3747_o_0),
    .Y(n_3957_o_0));
 OAI31xp33_ASAP7_75t_R n_3958 (.A1(net94),
    .A2(n_3684_o_0),
    .A3(n_3935_o_0),
    .B(n_3901_o_0),
    .Y(n_3958_o_0));
 AOI21xp33_ASAP7_75t_R n_3959 (.A1(n_3702_o_0),
    .A2(n_3958_o_0),
    .B(n_3748_o_0),
    .Y(n_3959_o_0));
 AOI31xp33_ASAP7_75t_R n_3960 (.A1(n_3627_o_0),
    .A2(n_3806_o_0),
    .A3(n_3766_o_0),
    .B(n_3702_o_0),
    .Y(n_3960_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3961 (.A1(n_3642_o_0),
    .A2(n_3739_o_0),
    .B(n_3755_o_0),
    .C(n_3960_o_0),
    .Y(n_3961_o_0));
 AOI22xp33_ASAP7_75t_R n_3962 (.A1(n_3954_o_0),
    .A2(n_3957_o_0),
    .B1(n_3959_o_0),
    .B2(n_3961_o_0),
    .Y(n_3962_o_0));
 INVx1_ASAP7_75t_R n_3963 (.A(n_3680_o_0),
    .Y(n_3963_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3964 (.A1(n_3801_o_0),
    .A2(n_3858_o_0),
    .B(n_3624_o_0),
    .C(n_3963_o_0),
    .Y(n_3964_o_0));
 NOR2xp33_ASAP7_75t_R n_3965 (.A(n_3659_o_0),
    .B(n_3683_o_0),
    .Y(n_3965_o_0));
 OAI21xp33_ASAP7_75t_R n_3966 (.A1(net74),
    .A2(n_3685_o_0),
    .B(n_3683_o_0),
    .Y(n_3966_o_0));
 NAND3xp33_ASAP7_75t_R n_3967 (.A(n_3750_o_0),
    .B(n_3966_o_0),
    .C(n_3627_o_0),
    .Y(n_3967_o_0));
 OAI31xp33_ASAP7_75t_R n_3968 (.A1(net11),
    .A2(n_3893_o_0),
    .A3(n_3965_o_0),
    .B(n_3967_o_0),
    .Y(n_3968_o_0));
 AOI21xp33_ASAP7_75t_R n_3969 (.A1(n_3700_o_0),
    .A2(n_3968_o_0),
    .B(n_3724_o_0),
    .Y(n_3969_o_0));
 AOI21xp33_ASAP7_75t_R n_3970 (.A1(n_3735_o_0),
    .A2(n_3732_o_0),
    .B(n_3705_o_0),
    .Y(n_3970_o_0));
 NAND2xp33_ASAP7_75t_R n_3971 (.A(n_3683_o_0),
    .B(n_3660_o_0),
    .Y(n_3971_o_0));
 OAI211xp5_ASAP7_75t_R n_3972 (.A1(net25),
    .A2(net72),
    .B(n_3971_o_0),
    .C(n_3627_o_0),
    .Y(n_3972_o_0));
 OAI211xp5_ASAP7_75t_R n_3973 (.A1(net11),
    .A2(n_3970_o_0),
    .B(n_3972_o_0),
    .C(n_3756_o_0),
    .Y(n_3973_o_0));
 INVx1_ASAP7_75t_R n_3974 (.A(n_3971_o_0),
    .Y(n_3974_o_0));
 AOI21xp33_ASAP7_75t_R n_3975 (.A1(n_3858_o_0),
    .A2(n_3800_o_0),
    .B(n_3700_o_0),
    .Y(n_3975_o_0));
 OAI31xp33_ASAP7_75t_R n_3976 (.A1(net11),
    .A2(n_3736_o_0),
    .A3(n_3974_o_0),
    .B(n_3975_o_0),
    .Y(n_3976_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3977 (.A1(n_3973_o_0),
    .A2(n_3976_o_0),
    .B(n_3748_o_0),
    .C(n_3604_o_0),
    .Y(n_3977_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_3978 (.A1(n_3756_o_0),
    .A2(n_3964_o_0),
    .B(n_3969_o_0),
    .C(n_3977_o_0),
    .Y(n_3978_o_0));
 AOI21xp33_ASAP7_75t_R n_3979 (.A1(n_3846_o_0),
    .A2(n_3962_o_0),
    .B(n_3978_o_0),
    .Y(n_3979_o_0));
 AOI21xp33_ASAP7_75t_R n_3980 (.A1(n_3821_o_0),
    .A2(n_3815_o_0),
    .B(n_3702_o_0),
    .Y(n_3980_o_0));
 OAI21xp33_ASAP7_75t_R n_3981 (.A1(n_3814_o_0),
    .A2(net11),
    .B(n_3980_o_0),
    .Y(n_3981_o_0));
 NAND2xp33_ASAP7_75t_R n_3982 (.A(n_3627_o_0),
    .B(n_3686_o_0),
    .Y(n_3982_o_0));
 AOI21xp33_ASAP7_75t_R n_3983 (.A1(n_3941_o_0),
    .A2(n_3882_o_0),
    .B(n_3700_o_0),
    .Y(n_3983_o_0));
 OAI21xp33_ASAP7_75t_R n_3984 (.A1(n_3982_o_0),
    .A2(n_3736_o_0),
    .B(n_3983_o_0),
    .Y(n_3984_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_3985 (.A1(n_3820_o_0),
    .A2(n_3859_o_0),
    .B(n_3981_o_0),
    .C(n_3984_o_0),
    .Y(n_3985_o_0));
 AO32x1_ASAP7_75t_R n_3986 (.A1(n_3712_o_0),
    .A2(n_3815_o_0),
    .A3(n_3627_o_0),
    .B1(n_3966_o_0),
    .B2(n_3941_o_0),
    .Y(n_3986_o_0));
 AOI21xp33_ASAP7_75t_R n_3987 (.A1(n_3770_o_0),
    .A2(n_3986_o_0),
    .B(n_3919_o_0),
    .Y(n_3987_o_0));
 OAI22xp33_ASAP7_75t_R n_3988 (.A1(n_3985_o_0),
    .A2(n_3723_o_0),
    .B1(n_3987_o_0),
    .B2(n_3747_o_0),
    .Y(n_3988_o_0));
 OAI21xp33_ASAP7_75t_R n_3989 (.A1(n_3798_o_0),
    .A2(n_3872_o_0),
    .B(n_3770_o_0),
    .Y(n_3989_o_0));
 OAI211xp5_ASAP7_75t_R n_3990 (.A1(n_3743_o_0),
    .A2(n_3790_o_0),
    .B(n_3776_o_0),
    .C(n_3627_o_0),
    .Y(n_3990_o_0));
 OAI21xp33_ASAP7_75t_R n_3991 (.A1(n_3912_o_0),
    .A2(n_3687_o_0),
    .B(net90),
    .Y(n_3991_o_0));
 AOI31xp33_ASAP7_75t_R n_3992 (.A1(n_3990_o_0),
    .A2(n_3991_o_0),
    .A3(n_3756_o_0),
    .B(n_3747_o_0),
    .Y(n_3992_o_0));
 OAI21xp33_ASAP7_75t_R n_3993 (.A1(n_3989_o_0),
    .A2(n_3767_o_0),
    .B(n_3992_o_0),
    .Y(n_3993_o_0));
 NAND3xp33_ASAP7_75t_R n_3994 (.A(n_3738_o_0),
    .B(n_3642_o_0),
    .C(net41),
    .Y(n_3994_o_0));
 NAND2xp33_ASAP7_75t_R n_3995 (.A(net93),
    .B(n_3736_o_0),
    .Y(n_3995_o_0));
 AOI21xp33_ASAP7_75t_R n_3996 (.A1(n_3994_o_0),
    .A2(n_3995_o_0),
    .B(n_3702_o_0),
    .Y(n_3996_o_0));
 OA21x2_ASAP7_75t_R n_3997 (.A1(net63),
    .A2(n_3912_o_0),
    .B(n_3915_o_0),
    .Y(n_3997_o_0));
 OAI21xp33_ASAP7_75t_R n_3998 (.A1(n_3996_o_0),
    .A2(n_3997_o_0),
    .B(n_3747_o_0),
    .Y(n_3998_o_0));
 AOI31xp33_ASAP7_75t_R n_3999 (.A1(n_3605_o_0),
    .A2(n_3993_o_0),
    .A3(n_3998_o_0),
    .B(n_3782_o_0),
    .Y(n_3999_o_0));
 OAI21xp33_ASAP7_75t_R n_4000 (.A1(n_3846_o_0),
    .A2(n_3988_o_0),
    .B(n_3999_o_0),
    .Y(n_4000_o_0));
 OAI21xp33_ASAP7_75t_R n_4001 (.A1(n_3613_o_0),
    .A2(n_3979_o_0),
    .B(n_4000_o_0),
    .Y(n_4001_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4002 (.A1(net25),
    .A2(net30),
    .B(n_3676_o_0),
    .C(net90),
    .Y(n_4002_o_0));
 AO21x1_ASAP7_75t_R n_4003 (.A1(n_3624_o_0),
    .A2(n_3805_o_0),
    .B(n_4002_o_0),
    .Y(n_4003_o_0));
 INVx1_ASAP7_75t_R n_4004 (.A(n_3780_o_0),
    .Y(n_4004_o_0));
 NOR4xp25_ASAP7_75t_R n_4005 (.A(n_3769_o_0),
    .B(n_3794_o_0),
    .C(n_3756_o_0),
    .D(net41),
    .Y(n_4005_o_0));
 AOI211xp5_ASAP7_75t_R n_4006 (.A1(n_3700_o_0),
    .A2(n_4003_o_0),
    .B(n_4004_o_0),
    .C(n_4005_o_0),
    .Y(n_4006_o_0));
 AOI211xp5_ASAP7_75t_R n_4007 (.A1(n_3660_o_0),
    .A2(net72),
    .B(n_3794_o_0),
    .C(net63),
    .Y(n_4007_o_0));
 AOI21xp33_ASAP7_75t_R n_4008 (.A1(n_3765_o_0),
    .A2(n_3971_o_0),
    .B(n_3624_o_0),
    .Y(n_4008_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4009 (.A1(n_3627_o_0),
    .A2(n_3685_o_0),
    .B(net72),
    .C(n_3702_o_0),
    .Y(n_4009_o_0));
 AOI21xp33_ASAP7_75t_R n_4010 (.A1(net63),
    .A2(n_3893_o_0),
    .B(n_4009_o_0),
    .Y(n_4010_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4011 (.A1(n_4007_o_0),
    .A2(n_4008_o_0),
    .B(n_3756_o_0),
    .C(n_4010_o_0),
    .Y(n_4011_o_0));
 AOI22xp33_ASAP7_75t_R n_4012 (.A1(n_4006_o_0),
    .A2(n_3605_o_0),
    .B1(n_3828_o_0),
    .B2(n_4011_o_0),
    .Y(n_4012_o_0));
 NAND3xp33_ASAP7_75t_R n_4013 (.A(n_3661_o_0),
    .B(n_3855_o_0),
    .C(n_3627_o_0),
    .Y(n_4013_o_0));
 OAI311xp33_ASAP7_75t_R n_4014 (.A1(net94),
    .A2(n_3939_o_0),
    .A3(n_3786_o_0),
    .B1(n_4013_o_0),
    .C1(n_3756_o_0),
    .Y(n_4014_o_0));
 INVx1_ASAP7_75t_R n_4015 (.A(n_3858_o_0),
    .Y(n_4015_o_0));
 OAI211xp5_ASAP7_75t_R n_4016 (.A1(n_3739_o_0),
    .A2(n_3705_o_0),
    .B(n_3627_o_0),
    .C(n_3710_o_0),
    .Y(n_4016_o_0));
 OAI31xp33_ASAP7_75t_R n_4017 (.A1(net94),
    .A2(n_3878_o_0),
    .A3(n_4015_o_0),
    .B(n_4016_o_0),
    .Y(n_4017_o_0));
 AOI21xp33_ASAP7_75t_R n_4018 (.A1(n_3702_o_0),
    .A2(n_4017_o_0),
    .B(n_3846_o_0),
    .Y(n_4018_o_0));
 NAND2xp33_ASAP7_75t_R n_4019 (.A(net90),
    .B(n_3811_o_0),
    .Y(n_4019_o_0));
 OAI22xp33_ASAP7_75t_R n_4020 (.A1(n_4019_o_0),
    .A2(n_3965_o_0),
    .B1(n_3810_o_0),
    .B2(n_4015_o_0),
    .Y(n_4020_o_0));
 OAI21xp33_ASAP7_75t_R n_4021 (.A1(n_3789_o_0),
    .A2(n_3624_o_0),
    .B(n_3702_o_0),
    .Y(n_4021_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4022 (.A1(net41),
    .A2(n_3769_o_0),
    .B(n_4021_o_0),
    .C(n_3605_o_0),
    .Y(n_4022_o_0));
 AOI21xp33_ASAP7_75t_R n_4023 (.A1(n_3700_o_0),
    .A2(n_4020_o_0),
    .B(n_4022_o_0),
    .Y(n_4023_o_0));
 AOI21xp33_ASAP7_75t_R n_4024 (.A1(n_4014_o_0),
    .A2(n_4018_o_0),
    .B(n_4023_o_0),
    .Y(n_4024_o_0));
 AOI22xp33_ASAP7_75t_R n_4025 (.A1(n_4012_o_0),
    .A2(n_3748_o_0),
    .B1(n_3724_o_0),
    .B2(n_4024_o_0),
    .Y(n_4025_o_0));
 NOR3xp33_ASAP7_75t_R n_4026 (.A(n_3737_o_0),
    .B(n_3965_o_0),
    .C(net11),
    .Y(n_4026_o_0));
 NAND3xp33_ASAP7_75t_R n_4027 (.A(n_3661_o_0),
    .B(n_3855_o_0),
    .C(n_3627_o_0),
    .Y(n_4027_o_0));
 INVx1_ASAP7_75t_R n_4028 (.A(n_4027_o_0),
    .Y(n_4028_o_0));
 OAI21xp33_ASAP7_75t_R n_4029 (.A1(n_4026_o_0),
    .A2(n_4028_o_0),
    .B(n_3700_o_0),
    .Y(n_4029_o_0));
 AO21x1_ASAP7_75t_R n_4030 (.A1(n_3679_o_0),
    .A2(n_3800_o_0),
    .B(n_3924_o_0),
    .Y(n_4030_o_0));
 AOI21xp33_ASAP7_75t_R n_4031 (.A1(n_3702_o_0),
    .A2(n_4030_o_0),
    .B(n_3846_o_0),
    .Y(n_4031_o_0));
 AOI21xp33_ASAP7_75t_R n_4032 (.A1(n_3814_o_0),
    .A2(n_4019_o_0),
    .B(n_3770_o_0),
    .Y(n_4032_o_0));
 NAND2xp33_ASAP7_75t_R n_4033 (.A(n_3702_o_0),
    .B(n_3787_o_0),
    .Y(n_4033_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4034 (.A1(net94),
    .A2(n_3708_o_0),
    .B(n_3824_o_0),
    .C(n_4033_o_0),
    .Y(n_4034_o_0));
 NOR3xp33_ASAP7_75t_R n_4035 (.A(n_4032_o_0),
    .B(n_4034_o_0),
    .C(n_3604_o_0),
    .Y(n_4035_o_0));
 AOI21xp33_ASAP7_75t_R n_4036 (.A1(n_4029_o_0),
    .A2(n_4031_o_0),
    .B(n_4035_o_0),
    .Y(n_4036_o_0));
 INVx1_ASAP7_75t_R n_4037 (.A(n_3912_o_0),
    .Y(n_4037_o_0));
 OAI21xp33_ASAP7_75t_R n_4038 (.A1(n_3627_o_0),
    .A2(n_3926_o_0),
    .B(n_4037_o_0),
    .Y(n_4038_o_0));
 INVx1_ASAP7_75t_R n_4039 (.A(n_3875_o_0),
    .Y(n_4039_o_0));
 INVx1_ASAP7_75t_R n_4040 (.A(n_3761_o_0),
    .Y(n_4040_o_0));
 NOR2xp33_ASAP7_75t_R n_4041 (.A(n_3626_o_0),
    .B(n_3684_o_0),
    .Y(n_4041_o_0));
 INVx1_ASAP7_75t_R n_4042 (.A(n_3970_o_0),
    .Y(n_4042_o_0));
 AOI21xp33_ASAP7_75t_R n_4043 (.A1(n_4041_o_0),
    .A2(n_4042_o_0),
    .B(n_3700_o_0),
    .Y(n_4043_o_0));
 OAI21xp33_ASAP7_75t_R n_4044 (.A1(n_4019_o_0),
    .A2(n_4040_o_0),
    .B(n_4043_o_0),
    .Y(n_4044_o_0));
 OAI311xp33_ASAP7_75t_R n_4045 (.A1(n_3702_o_0),
    .A2(n_4038_o_0),
    .A3(n_4039_o_0),
    .B1(n_3846_o_0),
    .C1(n_4044_o_0),
    .Y(n_4045_o_0));
 OAI22xp33_ASAP7_75t_R n_4046 (.A1(n_3879_o_0),
    .A2(n_3893_o_0),
    .B1(n_4040_o_0),
    .B2(n_3844_o_0),
    .Y(n_4046_o_0));
 AO21x1_ASAP7_75t_R n_4047 (.A1(n_3765_o_0),
    .A2(n_3679_o_0),
    .B(n_3627_o_0),
    .Y(n_4047_o_0));
 AOI31xp33_ASAP7_75t_R n_4048 (.A1(n_3770_o_0),
    .A2(n_3763_o_0),
    .A3(n_4047_o_0),
    .B(n_3605_o_0),
    .Y(n_4048_o_0));
 OAI21xp33_ASAP7_75t_R n_4049 (.A1(n_3702_o_0),
    .A2(n_4046_o_0),
    .B(n_4048_o_0),
    .Y(n_4049_o_0));
 AOI31xp33_ASAP7_75t_R n_4050 (.A1(n_3747_o_0),
    .A2(n_4045_o_0),
    .A3(n_4049_o_0),
    .B(n_3613_o_0),
    .Y(n_4050_o_0));
 OAI21xp33_ASAP7_75t_R n_4051 (.A1(n_3724_o_0),
    .A2(n_4036_o_0),
    .B(n_4050_o_0),
    .Y(n_4051_o_0));
 OAI21xp33_ASAP7_75t_R n_4052 (.A1(n_3782_o_0),
    .A2(n_4025_o_0),
    .B(n_4051_o_0),
    .Y(n_4052_o_0));
 INVx1_ASAP7_75t_R n_4053 (.A(n_3982_o_0),
    .Y(n_4053_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4054 (.A1(n_3815_o_0),
    .A2(n_3712_o_0),
    .B(net11),
    .C(n_3756_o_0),
    .Y(n_4054_o_0));
 AOI21xp33_ASAP7_75t_R n_4055 (.A1(n_3855_o_0),
    .A2(n_4053_o_0),
    .B(n_4054_o_0),
    .Y(n_4055_o_0));
 AOI21xp33_ASAP7_75t_R n_4056 (.A1(n_3907_o_0),
    .A2(n_4027_o_0),
    .B(n_3756_o_0),
    .Y(n_4056_o_0));
 AOI32xp33_ASAP7_75t_R n_4057 (.A1(n_3894_o_0),
    .A2(n_4002_o_0),
    .A3(n_3756_o_0),
    .B1(n_3769_o_0),
    .B2(net90),
    .Y(n_4057_o_0));
 NOR4xp25_ASAP7_75t_R n_4058 (.A(n_3820_o_0),
    .B(n_3756_o_0),
    .C(n_3627_o_0),
    .D(n_3705_o_0),
    .Y(n_4058_o_0));
 NOR2xp33_ASAP7_75t_R n_4059 (.A(n_3642_o_0),
    .B(n_3738_o_0),
    .Y(n_4059_o_0));
 OAI31xp33_ASAP7_75t_R n_4060 (.A1(net63),
    .A2(n_4059_o_0),
    .A3(n_3736_o_0),
    .B(n_3911_o_0),
    .Y(n_4060_o_0));
 OAI221xp5_ASAP7_75t_R n_4061 (.A1(n_4057_o_0),
    .A2(n_4058_o_0),
    .B1(n_3700_o_0),
    .B2(n_4060_o_0),
    .C(n_3604_o_0),
    .Y(n_4061_o_0));
 OAI31xp33_ASAP7_75t_R n_4062 (.A1(n_3828_o_0),
    .A2(n_4055_o_0),
    .A3(n_4056_o_0),
    .B(n_4061_o_0),
    .Y(n_4062_o_0));
 OA21x2_ASAP7_75t_R n_4063 (.A1(n_3721_o_0),
    .A2(n_3722_o_0),
    .B(n_4062_o_0),
    .Y(n_4063_o_0));
 NOR2xp33_ASAP7_75t_R n_4064 (.A(n_3756_o_0),
    .B(n_3804_o_0),
    .Y(n_4064_o_0));
 AOI21xp33_ASAP7_75t_R n_4065 (.A1(n_3858_o_0),
    .A2(n_3859_o_0),
    .B(n_3702_o_0),
    .Y(n_4065_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4066 (.A1(net41),
    .A2(n_3794_o_0),
    .B(n_4065_o_0),
    .C(n_3605_o_0),
    .Y(n_4066_o_0));
 INVx1_ASAP7_75t_R n_4067 (.A(n_4066_o_0),
    .Y(n_4067_o_0));
 AOI21xp33_ASAP7_75t_R n_4068 (.A1(n_3991_o_0),
    .A2(n_4064_o_0),
    .B(n_4067_o_0),
    .Y(n_4068_o_0));
 AOI211xp5_ASAP7_75t_R n_4069 (.A1(net30),
    .A2(n_3786_o_0),
    .B(n_3744_o_0),
    .C(n_3624_o_0),
    .Y(n_4069_o_0));
 AOI31xp33_ASAP7_75t_R n_4070 (.A1(n_3624_o_0),
    .A2(n_3685_o_0),
    .A3(n_3762_o_0),
    .B(n_4069_o_0),
    .Y(n_4070_o_0));
 AOI21xp33_ASAP7_75t_R n_4071 (.A1(net25),
    .A2(net30),
    .B(n_3743_o_0),
    .Y(n_4071_o_0));
 OAI31xp33_ASAP7_75t_R n_4072 (.A1(n_3627_o_0),
    .A2(n_3794_o_0),
    .A3(n_4071_o_0),
    .B(n_3770_o_0),
    .Y(n_4072_o_0));
 AOI31xp33_ASAP7_75t_R n_4073 (.A1(n_3679_o_0),
    .A2(n_3627_o_0),
    .A3(n_3710_o_0),
    .B(n_4072_o_0),
    .Y(n_4073_o_0));
 AOI211xp5_ASAP7_75t_R n_4074 (.A1(n_3756_o_0),
    .A2(n_4070_o_0),
    .B(n_4073_o_0),
    .C(n_3828_o_0),
    .Y(n_4074_o_0));
 NOR3xp33_ASAP7_75t_R n_4075 (.A(n_4068_o_0),
    .B(n_4074_o_0),
    .C(n_3724_o_0),
    .Y(n_4075_o_0));
 AO21x1_ASAP7_75t_R n_4076 (.A1(n_3875_o_0),
    .A2(n_3791_o_0),
    .B(n_3828_o_0),
    .Y(n_4076_o_0));
 INVx1_ASAP7_75t_R n_4077 (.A(n_3750_o_0),
    .Y(n_4077_o_0));
 OAI311xp33_ASAP7_75t_R n_4078 (.A1(n_3685_o_0),
    .A2(n_3705_o_0),
    .A3(net30),
    .B1(n_3624_o_0),
    .C1(n_3776_o_0),
    .Y(n_4078_o_0));
 OAI31xp33_ASAP7_75t_R n_4079 (.A1(net41),
    .A2(n_3893_o_0),
    .A3(n_4077_o_0),
    .B(n_4078_o_0),
    .Y(n_4079_o_0));
 AOI21xp33_ASAP7_75t_R n_4080 (.A1(n_3604_o_0),
    .A2(n_4079_o_0),
    .B(n_3702_o_0),
    .Y(n_4080_o_0));
 OAI21xp33_ASAP7_75t_R n_4081 (.A1(net30),
    .A2(n_3685_o_0),
    .B(n_3624_o_0),
    .Y(n_4081_o_0));
 OAI21xp33_ASAP7_75t_R n_4082 (.A1(net41),
    .A2(n_3940_o_0),
    .B(n_4081_o_0),
    .Y(n_4082_o_0));
 AOI21xp33_ASAP7_75t_R n_4083 (.A1(n_3941_o_0),
    .A2(n_3846_o_0),
    .B(n_3700_o_0),
    .Y(n_4083_o_0));
 OAI21xp33_ASAP7_75t_R n_4084 (.A1(n_3940_o_0),
    .A2(n_3945_o_0),
    .B(n_4083_o_0),
    .Y(n_4084_o_0));
 AOI21xp33_ASAP7_75t_R n_4085 (.A1(n_3604_o_0),
    .A2(n_4082_o_0),
    .B(n_4084_o_0),
    .Y(n_4085_o_0));
 AOI21xp33_ASAP7_75t_R n_4086 (.A1(n_4076_o_0),
    .A2(n_4080_o_0),
    .B(n_4085_o_0),
    .Y(n_4086_o_0));
 AOI21xp33_ASAP7_75t_R n_4087 (.A1(n_3744_o_0),
    .A2(n_3624_o_0),
    .B(n_3846_o_0),
    .Y(n_4087_o_0));
 NAND3xp33_ASAP7_75t_R n_4088 (.A(n_3882_o_0),
    .B(n_3712_o_0),
    .C(n_3627_o_0),
    .Y(n_4088_o_0));
 OAI31xp33_ASAP7_75t_R n_4089 (.A1(n_3624_o_0),
    .A2(n_3965_o_0),
    .A3(n_3744_o_0),
    .B(n_3605_o_0),
    .Y(n_4089_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4090 (.A1(n_3963_o_0),
    .A2(n_3832_o_0),
    .B(n_4089_o_0),
    .C(n_3700_o_0),
    .Y(n_4090_o_0));
 AO21x1_ASAP7_75t_R n_4091 (.A1(net25),
    .A2(n_3624_o_0),
    .B(n_3800_o_0),
    .Y(n_4091_o_0));
 AOI32xp33_ASAP7_75t_R n_4092 (.A1(n_3624_o_0),
    .A2(n_3712_o_0),
    .A3(n_3686_o_0),
    .B1(net25),
    .B2(n_3742_o_0),
    .Y(n_4092_o_0));
 AOI31xp33_ASAP7_75t_R n_4093 (.A1(n_3875_o_0),
    .A2(n_4092_o_0),
    .A3(n_3828_o_0),
    .B(n_3756_o_0),
    .Y(n_4093_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4094 (.A1(n_3799_o_0),
    .A2(n_4091_o_0),
    .B(n_3604_o_0),
    .C(n_4093_o_0),
    .Y(n_4094_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4095 (.A1(n_4087_o_0),
    .A2(n_4088_o_0),
    .B(n_4090_o_0),
    .C(n_4094_o_0),
    .Y(n_4095_o_0));
 OAI221xp5_ASAP7_75t_R n_4096 (.A1(n_3748_o_0),
    .A2(n_4086_o_0),
    .B1(n_3724_o_0),
    .B2(n_4095_o_0),
    .C(n_3613_o_0),
    .Y(n_4096_o_0));
 OAI31xp33_ASAP7_75t_R n_4097 (.A1(n_4063_o_0),
    .A2(n_4075_o_0),
    .A3(n_3613_o_0),
    .B(n_4096_o_0),
    .Y(n_4097_o_0));
 NOR3xp33_ASAP7_75t_R n_4098 (.A(n_3709_o_0),
    .B(n_3682_o_0),
    .C(net25),
    .Y(n_4098_o_0));
 OAI31xp33_ASAP7_75t_R n_4099 (.A1(n_3774_o_0),
    .A2(n_4098_o_0),
    .A3(n_3627_o_0),
    .B(n_3771_o_0),
    .Y(n_4099_o_0));
 AOI21xp33_ASAP7_75t_R n_4100 (.A1(net94),
    .A2(n_3900_o_0),
    .B(n_4099_o_0),
    .Y(n_4100_o_0));
 NOR3xp33_ASAP7_75t_R n_4101 (.A(n_3744_o_0),
    .B(n_3624_o_0),
    .C(n_3684_o_0),
    .Y(n_4101_o_0));
 AOI31xp33_ASAP7_75t_R n_4102 (.A1(n_3624_o_0),
    .A2(n_3710_o_0),
    .A3(n_3805_o_0),
    .B(n_4101_o_0),
    .Y(n_4102_o_0));
 NOR2xp33_ASAP7_75t_R n_4103 (.A(n_3756_o_0),
    .B(n_4102_o_0),
    .Y(n_4103_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4104 (.A1(n_3660_o_0),
    .A2(net94),
    .B(n_3843_o_0),
    .C(n_3858_o_0),
    .Y(n_4104_o_0));
 OAI31xp33_ASAP7_75t_R n_4105 (.A1(net63),
    .A2(n_3739_o_0),
    .A3(n_3642_o_0),
    .B(n_3937_o_0),
    .Y(n_4105_o_0));
 AO21x1_ASAP7_75t_R n_4106 (.A1(n_3774_o_0),
    .A2(n_3624_o_0),
    .B(n_4105_o_0),
    .Y(n_4106_o_0));
 AOI21xp33_ASAP7_75t_R n_4107 (.A1(n_3700_o_0),
    .A2(n_4106_o_0),
    .B(n_3604_o_0),
    .Y(n_4107_o_0));
 OAI21xp33_ASAP7_75t_R n_4108 (.A1(n_3756_o_0),
    .A2(n_4104_o_0),
    .B(n_4107_o_0),
    .Y(n_4108_o_0));
 OAI311xp33_ASAP7_75t_R n_4109 (.A1(n_3846_o_0),
    .A2(n_4100_o_0),
    .A3(n_4103_o_0),
    .B1(n_3748_o_0),
    .C1(n_4108_o_0),
    .Y(n_4109_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4110 (.A1(n_3682_o_0),
    .A2(n_3709_o_0),
    .B(net25),
    .C(n_3867_o_0),
    .Y(n_4110_o_0));
 AOI31xp33_ASAP7_75t_R n_4111 (.A1(n_3624_o_0),
    .A2(n_3761_o_0),
    .A3(n_3766_o_0),
    .B(n_4110_o_0),
    .Y(n_4111_o_0));
 OAI211xp5_ASAP7_75t_R n_4112 (.A1(n_3705_o_0),
    .A2(n_3738_o_0),
    .B(n_3750_o_0),
    .C(n_3627_o_0),
    .Y(n_4112_o_0));
 OAI31xp33_ASAP7_75t_R n_4113 (.A1(net94),
    .A2(n_3680_o_0),
    .A3(n_3965_o_0),
    .B(n_4112_o_0),
    .Y(n_4113_o_0));
 AOI21xp33_ASAP7_75t_R n_4114 (.A1(n_3846_o_0),
    .A2(n_4113_o_0),
    .B(n_3700_o_0),
    .Y(n_4114_o_0));
 OAI21xp33_ASAP7_75t_R n_4115 (.A1(n_3605_o_0),
    .A2(n_4111_o_0),
    .B(n_4114_o_0),
    .Y(n_4115_o_0));
 NAND2xp33_ASAP7_75t_R n_4116 (.A(n_3995_o_0),
    .B(n_3946_o_0),
    .Y(n_4116_o_0));
 NOR3xp33_ASAP7_75t_R n_4117 (.A(n_4015_o_0),
    .B(n_3708_o_0),
    .C(net63),
    .Y(n_4117_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4118 (.A1(n_3744_o_0),
    .A2(n_3627_o_0),
    .B(n_4117_o_0),
    .C(n_3604_o_0),
    .Y(n_4118_o_0));
 OAI211xp5_ASAP7_75t_R n_4119 (.A1(n_4116_o_0),
    .A2(n_3828_o_0),
    .B(n_4118_o_0),
    .C(n_3756_o_0),
    .Y(n_4119_o_0));
 AOI31xp33_ASAP7_75t_R n_4120 (.A1(n_3724_o_0),
    .A2(n_4115_o_0),
    .A3(n_4119_o_0),
    .B(n_3613_o_0),
    .Y(n_4120_o_0));
 NOR2xp33_ASAP7_75t_R n_4121 (.A(net93),
    .B(n_3708_o_0),
    .Y(n_4121_o_0));
 AOI21xp33_ASAP7_75t_R n_4122 (.A1(n_3787_o_0),
    .A2(n_3788_o_0),
    .B(n_4121_o_0),
    .Y(n_4122_o_0));
 AOI31xp33_ASAP7_75t_R n_4123 (.A1(n_3624_o_0),
    .A2(n_4037_o_0),
    .A3(n_3686_o_0),
    .B(n_3700_o_0),
    .Y(n_4123_o_0));
 AOI21xp33_ASAP7_75t_R n_4124 (.A1(n_3751_o_0),
    .A2(n_4123_o_0),
    .B(n_3846_o_0),
    .Y(n_4124_o_0));
 NAND2xp33_ASAP7_75t_R n_4125 (.A(n_3766_o_0),
    .B(n_3700_o_0),
    .Y(n_4125_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4126 (.A1(net11),
    .A2(n_3798_o_0),
    .B(n_3835_o_0),
    .C(n_4125_o_0),
    .Y(n_4126_o_0));
 OAI21xp33_ASAP7_75t_R n_4127 (.A1(n_3685_o_0),
    .A2(net93),
    .B(n_3660_o_0),
    .Y(n_4127_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4128 (.A1(n_3685_o_0),
    .A2(n_3642_o_0),
    .B(n_4127_o_0),
    .C(n_3756_o_0),
    .Y(n_4128_o_0));
 NOR3xp33_ASAP7_75t_R n_4129 (.A(n_4126_o_0),
    .B(n_4128_o_0),
    .C(n_3604_o_0),
    .Y(n_4129_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4130 (.A1(n_3770_o_0),
    .A2(n_4122_o_0),
    .B(n_4124_o_0),
    .C(n_4129_o_0),
    .Y(n_4130_o_0));
 NOR3xp33_ASAP7_75t_R n_4131 (.A(n_3744_o_0),
    .B(n_3627_o_0),
    .C(n_3965_o_0),
    .Y(n_4131_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4132 (.A1(n_3627_o_0),
    .A2(n_3815_o_0),
    .B(n_4131_o_0),
    .C(n_3700_o_0),
    .Y(n_4132_o_0));
 OA21x2_ASAP7_75t_R n_4133 (.A1(n_3898_o_0),
    .A2(n_3756_o_0),
    .B(n_3828_o_0),
    .Y(n_4133_o_0));
 NAND2xp33_ASAP7_75t_R n_4134 (.A(net30),
    .B(n_3683_o_0),
    .Y(n_4134_o_0));
 OAI21xp33_ASAP7_75t_R n_4135 (.A1(net72),
    .A2(net30),
    .B(n_4134_o_0),
    .Y(n_4135_o_0));
 INVx1_ASAP7_75t_R n_4136 (.A(n_4135_o_0),
    .Y(n_4136_o_0));
 AOI31xp33_ASAP7_75t_R n_4137 (.A1(net63),
    .A2(n_3811_o_0),
    .A3(n_3661_o_0),
    .B(n_3700_o_0),
    .Y(n_4137_o_0));
 OAI21xp33_ASAP7_75t_R n_4138 (.A1(net11),
    .A2(n_4136_o_0),
    .B(n_4137_o_0),
    .Y(n_4138_o_0));
 OAI31xp33_ASAP7_75t_R n_4139 (.A1(net94),
    .A2(n_3893_o_0),
    .A3(n_4077_o_0),
    .B(n_3840_o_0),
    .Y(n_4139_o_0));
 AOI21xp33_ASAP7_75t_R n_4140 (.A1(n_4138_o_0),
    .A2(n_4139_o_0),
    .B(n_3604_o_0),
    .Y(n_4140_o_0));
 AOI211xp5_ASAP7_75t_R n_4141 (.A1(n_4132_o_0),
    .A2(n_4133_o_0),
    .B(n_4140_o_0),
    .C(n_3723_o_0),
    .Y(n_4141_o_0));
 AOI211xp5_ASAP7_75t_R n_4142 (.A1(n_4130_o_0),
    .A2(n_3748_o_0),
    .B(n_4141_o_0),
    .C(n_3782_o_0),
    .Y(n_4142_o_0));
 AOI21xp33_ASAP7_75t_R n_4143 (.A1(n_4109_o_0),
    .A2(n_4120_o_0),
    .B(n_4142_o_0),
    .Y(n_4143_o_0));
 NAND2xp33_ASAP7_75t_R n_4144 (.A(n_3604_o_0),
    .B(n_3995_o_0),
    .Y(n_4144_o_0));
 AOI31xp33_ASAP7_75t_R n_4145 (.A1(n_3624_o_0),
    .A2(n_3799_o_0),
    .A3(n_3894_o_0),
    .B(n_3604_o_0),
    .Y(n_4145_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4146 (.A1(net25),
    .A2(n_3708_o_0),
    .B(n_3662_o_0),
    .C(n_4145_o_0),
    .Y(n_4146_o_0));
 OAI211xp5_ASAP7_75t_R n_4147 (.A1(n_4144_o_0),
    .A2(n_3857_o_0),
    .B(n_3702_o_0),
    .C(n_4146_o_0),
    .Y(n_4147_o_0));
 AOI22xp33_ASAP7_75t_R n_4148 (.A1(n_4121_o_0),
    .A2(n_3787_o_0),
    .B1(n_3627_o_0),
    .B2(n_3685_o_0),
    .Y(n_4148_o_0));
 AOI31xp33_ASAP7_75t_R n_4149 (.A1(n_3627_o_0),
    .A2(n_3750_o_0),
    .A3(n_3805_o_0),
    .B(n_3846_o_0),
    .Y(n_4149_o_0));
 OAI21xp33_ASAP7_75t_R n_4150 (.A1(net94),
    .A2(n_4040_o_0),
    .B(n_4149_o_0),
    .Y(n_4150_o_0));
 OAI211xp5_ASAP7_75t_R n_4151 (.A1(n_3604_o_0),
    .A2(n_4148_o_0),
    .B(n_4150_o_0),
    .C(n_3700_o_0),
    .Y(n_4151_o_0));
 AND3x1_ASAP7_75t_R n_4152 (.A(n_4147_o_0),
    .B(n_4151_o_0),
    .C(n_3747_o_0),
    .Y(n_4152_o_0));
 AOI21xp33_ASAP7_75t_R n_4153 (.A1(n_4041_o_0),
    .A2(n_3966_o_0),
    .B(n_3846_o_0),
    .Y(n_4153_o_0));
 NOR3xp33_ASAP7_75t_R n_4154 (.A(n_4131_o_0),
    .B(n_3604_o_0),
    .C(n_4041_o_0),
    .Y(n_4154_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4155 (.A1(n_3786_o_0),
    .A2(n_3844_o_0),
    .B(n_4153_o_0),
    .C(n_4154_o_0),
    .Y(n_4155_o_0));
 NAND3xp33_ASAP7_75t_R n_4156 (.A(n_3661_o_0),
    .B(n_3627_o_0),
    .C(n_3685_o_0),
    .Y(n_4156_o_0));
 AOI21xp33_ASAP7_75t_R n_4157 (.A1(n_3765_o_0),
    .A2(n_3971_o_0),
    .B(n_3627_o_0),
    .Y(n_4157_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4158 (.A1(net11),
    .A2(n_3687_o_0),
    .B(n_4156_o_0),
    .C(n_4157_o_0),
    .Y(n_4158_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4159 (.A1(n_3776_o_0),
    .A2(n_4053_o_0),
    .B(n_3871_o_0),
    .C(n_3700_o_0),
    .Y(n_4159_o_0));
 AOI21xp33_ASAP7_75t_R n_4160 (.A1(n_3605_o_0),
    .A2(n_4158_o_0),
    .B(n_4159_o_0),
    .Y(n_4160_o_0));
 AOI211xp5_ASAP7_75t_R n_4161 (.A1(n_3702_o_0),
    .A2(n_4155_o_0),
    .B(n_4160_o_0),
    .C(n_3724_o_0),
    .Y(n_4161_o_0));
 AOI21xp33_ASAP7_75t_R n_4162 (.A1(net30),
    .A2(n_3801_o_0),
    .B(n_3624_o_0),
    .Y(n_4162_o_0));
 OAI21xp33_ASAP7_75t_R n_4163 (.A1(net11),
    .A2(n_3790_o_0),
    .B(n_3759_o_0),
    .Y(n_4163_o_0));
 OAI31xp33_ASAP7_75t_R n_4164 (.A1(n_3770_o_0),
    .A2(n_4007_o_0),
    .A3(n_4162_o_0),
    .B(n_4163_o_0),
    .Y(n_4164_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4165 (.A1(n_3641_o_0),
    .A2(n_3637_o_0),
    .B(n_3820_o_0),
    .C(n_3754_o_0),
    .Y(n_4165_o_0));
 OAI31xp33_ASAP7_75t_R n_4166 (.A1(n_3965_o_0),
    .A2(n_3687_o_0),
    .A3(net41),
    .B(n_4165_o_0),
    .Y(n_4166_o_0));
 NOR3xp33_ASAP7_75t_R n_4167 (.A(n_4166_o_0),
    .B(n_3770_o_0),
    .C(n_3605_o_0),
    .Y(n_4167_o_0));
 OR2x2_ASAP7_75t_R n_4168 (.A(_00921_),
    .B(n_3602_o_0),
    .Y(n_4168_o_0));
 OAI21xp33_ASAP7_75t_R n_4169 (.A1(n_3912_o_0),
    .A2(n_3970_o_0),
    .B(net63),
    .Y(n_4169_o_0));
 OAI31xp33_ASAP7_75t_R n_4170 (.A1(n_3642_o_0),
    .A2(net30),
    .A3(n_3627_o_0),
    .B(n_4169_o_0),
    .Y(n_4170_o_0));
 AOI211xp5_ASAP7_75t_R n_4171 (.A1(n_4168_o_0),
    .A2(n_3603_o_0),
    .B(n_4170_o_0),
    .C(n_3700_o_0),
    .Y(n_4171_o_0));
 AOI211xp5_ASAP7_75t_R n_4172 (.A1(n_3846_o_0),
    .A2(n_4164_o_0),
    .B(n_4167_o_0),
    .C(n_4171_o_0),
    .Y(n_4172_o_0));
 AOI21xp33_ASAP7_75t_R n_4173 (.A1(n_3858_o_0),
    .A2(n_3843_o_0),
    .B(n_3702_o_0),
    .Y(n_4173_o_0));
 OAI21xp33_ASAP7_75t_R n_4174 (.A1(n_3779_o_0),
    .A2(net41),
    .B(n_4173_o_0),
    .Y(n_4174_o_0));
 OAI31xp33_ASAP7_75t_R n_4175 (.A1(n_3938_o_0),
    .A2(n_3760_o_0),
    .A3(n_4157_o_0),
    .B(n_4174_o_0),
    .Y(n_4175_o_0));
 AOI21xp33_ASAP7_75t_R n_4176 (.A1(n_3966_o_0),
    .A2(n_3941_o_0),
    .B(n_3702_o_0),
    .Y(n_4176_o_0));
 OAI21xp33_ASAP7_75t_R n_4177 (.A1(n_3872_o_0),
    .A2(n_3856_o_0),
    .B(n_4176_o_0),
    .Y(n_4177_o_0));
 AOI31xp33_ASAP7_75t_R n_4178 (.A1(n_3624_o_0),
    .A2(n_3750_o_0),
    .A3(n_3815_o_0),
    .B(n_3700_o_0),
    .Y(n_4178_o_0));
 AO31x2_ASAP7_75t_R n_4179 (.A1(n_3686_o_0),
    .A2(n_3765_o_0),
    .A3(n_3971_o_0),
    .B(n_3624_o_0),
    .Y(n_4179_o_0));
 AOI21xp33_ASAP7_75t_R n_4180 (.A1(n_4178_o_0),
    .A2(n_4179_o_0),
    .B(n_3828_o_0),
    .Y(n_4180_o_0));
 AOI21xp33_ASAP7_75t_R n_4181 (.A1(n_4177_o_0),
    .A2(n_4180_o_0),
    .B(n_3724_o_0),
    .Y(n_4181_o_0));
 OAI21xp33_ASAP7_75t_R n_4182 (.A1(n_3605_o_0),
    .A2(n_4175_o_0),
    .B(n_4181_o_0),
    .Y(n_4182_o_0));
 OAI211xp5_ASAP7_75t_R n_4183 (.A1(n_4172_o_0),
    .A2(n_3723_o_0),
    .B(n_4182_o_0),
    .C(n_3782_o_0),
    .Y(n_4183_o_0));
 OAI31xp33_ASAP7_75t_R n_4184 (.A1(n_3782_o_0),
    .A2(n_4152_o_0),
    .A3(n_4161_o_0),
    .B(n_4183_o_0),
    .Y(n_4184_o_0));
 XNOR2xp5_ASAP7_75t_R n_4185 (.A(_01013_),
    .B(_01053_),
    .Y(n_4185_o_0));
 XOR2xp5_ASAP7_75t_R n_4186 (.A(_01062_),
    .B(_01101_),
    .Y(n_4186_o_0));
 NAND2xp33_ASAP7_75t_R n_4187 (.A(_01054_),
    .B(n_4186_o_0),
    .Y(n_4187_o_0));
 OAI21xp33_ASAP7_75t_R n_4188 (.A1(_01054_),
    .A2(n_4186_o_0),
    .B(n_4187_o_0),
    .Y(n_4188_o_0));
 NOR2xp33_ASAP7_75t_R n_4189 (.A(n_4185_o_0),
    .B(n_4188_o_0),
    .Y(n_4189_o_0));
 AO21x1_ASAP7_75t_R n_4190 (.A1(n_4185_o_0),
    .A2(n_4188_o_0),
    .B(n_4189_o_0),
    .Y(n_4190_o_0));
 OAI21xp33_ASAP7_75t_R n_4191 (.A1(_00512_),
    .A2(net77),
    .B(n_2462_o_0),
    .Y(n_4191_o_0));
 INVx1_ASAP7_75t_R n_4192 (.A(_00512_),
    .Y(n_4192_o_0));
 AOI21xp33_ASAP7_75t_R n_4193 (.A1(n_4185_o_0),
    .A2(n_4188_o_0),
    .B(n_3021_o_0),
    .Y(n_4193_o_0));
 INVx1_ASAP7_75t_R n_4194 (.A(n_4185_o_0),
    .Y(n_4194_o_0));
 XNOR2xp5_ASAP7_75t_R n_4195 (.A(_01062_),
    .B(_01101_),
    .Y(n_4195_o_0));
 XNOR2xp5_ASAP7_75t_R n_4196 (.A(_01054_),
    .B(n_4195_o_0),
    .Y(n_4196_o_0));
 NAND2xp33_ASAP7_75t_R n_4197 (.A(n_4194_o_0),
    .B(n_4196_o_0),
    .Y(n_4197_o_0));
 AOI21xp33_ASAP7_75t_R n_4198 (.A1(n_4193_o_0),
    .A2(n_4197_o_0),
    .B(n_2462_o_0),
    .Y(n_4198_o_0));
 OAI21xp33_ASAP7_75t_R n_4199 (.A1(n_4192_o_0),
    .A2(net),
    .B(n_4198_o_0),
    .Y(n_4199_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4200 (.A1(n_4190_o_0),
    .A2(net),
    .B(n_4191_o_0),
    .C(n_4199_o_0),
    .Y(n_4200_o_0));
 XNOR2xp5_ASAP7_75t_R n_4201 (.A(_01012_),
    .B(_01019_),
    .Y(n_4201_o_0));
 INVx1_ASAP7_75t_R n_4202 (.A(_01100_),
    .Y(n_4202_o_0));
 NAND2xp33_ASAP7_75t_R n_4203 (.A(n_4202_o_0),
    .B(n_4201_o_0),
    .Y(n_4203_o_0));
 OAI21xp33_ASAP7_75t_R n_4204 (.A1(n_4201_o_0),
    .A2(n_4202_o_0),
    .B(n_4203_o_0),
    .Y(n_4204_o_0));
 XNOR2xp5_ASAP7_75t_R n_4205 (.A(_01052_),
    .B(_01059_),
    .Y(n_4205_o_0));
 XNOR2xp5_ASAP7_75t_R n_4206 (.A(_01053_),
    .B(_01061_),
    .Y(n_4206_o_0));
 NAND2xp33_ASAP7_75t_R n_4207 (.A(n_4206_o_0),
    .B(n_4205_o_0),
    .Y(n_4207_o_0));
 OAI21xp33_ASAP7_75t_R n_4208 (.A1(n_4205_o_0),
    .A2(n_4206_o_0),
    .B(n_4207_o_0),
    .Y(n_4208_o_0));
 XOR2xp5_ASAP7_75t_R n_4209 (.A(_01052_),
    .B(_01059_),
    .Y(n_4209_o_0));
 XOR2xp5_ASAP7_75t_R n_4210 (.A(_01053_),
    .B(_01061_),
    .Y(n_4210_o_0));
 NOR2xp33_ASAP7_75t_R n_4211 (.A(n_4209_o_0),
    .B(n_4210_o_0),
    .Y(n_4211_o_0));
 NOR2xp33_ASAP7_75t_R n_4212 (.A(n_4206_o_0),
    .B(n_4205_o_0),
    .Y(n_4212_o_0));
 XOR2xp5_ASAP7_75t_R n_4213 (.A(_01012_),
    .B(_01019_),
    .Y(n_4213_o_0));
 NOR2xp33_ASAP7_75t_R n_4214 (.A(_01100_),
    .B(n_4213_o_0),
    .Y(n_4214_o_0));
 NOR2xp33_ASAP7_75t_R n_4215 (.A(n_4202_o_0),
    .B(n_4201_o_0),
    .Y(n_4215_o_0));
 OAI22xp33_ASAP7_75t_R n_4216 (.A1(n_4211_o_0),
    .A2(n_4212_o_0),
    .B1(n_4214_o_0),
    .B2(n_4215_o_0),
    .Y(n_4216_o_0));
 OAI21xp33_ASAP7_75t_R n_4217 (.A1(n_4204_o_0),
    .A2(n_4208_o_0),
    .B(n_4216_o_0),
    .Y(n_4217_o_0));
 AOI21xp33_ASAP7_75t_R n_4218 (.A1(_00509_),
    .A2(net5),
    .B(n_2445_o_0),
    .Y(n_4218_o_0));
 XNOR2xp5_ASAP7_75t_R n_4219 (.A(_01100_),
    .B(n_4201_o_0),
    .Y(n_4219_o_0));
 XNOR2xp5_ASAP7_75t_R n_4220 (.A(n_4205_o_0),
    .B(n_4210_o_0),
    .Y(n_4220_o_0));
 NAND2xp33_ASAP7_75t_R n_4221 (.A(n_4209_o_0),
    .B(n_4210_o_0),
    .Y(n_4221_o_0));
 NAND2xp33_ASAP7_75t_R n_4222 (.A(_01100_),
    .B(n_4213_o_0),
    .Y(n_4222_o_0));
 AOI22xp33_ASAP7_75t_R n_4223 (.A1(n_4221_o_0),
    .A2(n_4207_o_0),
    .B1(n_4203_o_0),
    .B2(n_4222_o_0),
    .Y(n_4223_o_0));
 OAI21xp33_ASAP7_75t_R n_4224 (.A1(_00509_),
    .A2(_00858_),
    .B(n_2445_o_0),
    .Y(n_4224_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4225 (.A1(n_4219_o_0),
    .A2(n_4220_o_0),
    .B(n_4223_o_0),
    .C(net77),
    .D(n_4224_o_0),
    .Y(n_4225_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_4226 (.A1(n_3021_o_0),
    .A2(n_4217_o_0),
    .B(n_4218_o_0),
    .C(n_4225_o_0),
    .Y(n_4226_o_0));
 XNOR2xp5_ASAP7_75t_R n_4227 (.A(_01019_),
    .B(_01059_),
    .Y(n_4227_o_0));
 INVx1_ASAP7_75t_R n_4228 (.A(_01099_),
    .Y(n_4228_o_0));
 NAND2xp33_ASAP7_75t_R n_4229 (.A(n_4228_o_0),
    .B(n_4227_o_0),
    .Y(n_4229_o_0));
 XNOR2xp5_ASAP7_75t_R n_4230 (.A(_01052_),
    .B(_01060_),
    .Y(n_4230_o_0));
 INVx1_ASAP7_75t_R n_4231 (.A(n_4230_o_0),
    .Y(n_4231_o_0));
 OAI211xp5_ASAP7_75t_R n_4232 (.A1(n_4227_o_0),
    .A2(n_4228_o_0),
    .B(n_4229_o_0),
    .C(n_4231_o_0),
    .Y(n_4232_o_0));
 NOR2xp33_ASAP7_75t_R n_4233 (.A(n_4228_o_0),
    .B(n_4227_o_0),
    .Y(n_4233_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4234 (.A1(n_4227_o_0),
    .A2(n_4228_o_0),
    .B(n_4233_o_0),
    .C(n_4230_o_0),
    .Y(n_4234_o_0));
 NOR2xp33_ASAP7_75t_R n_4235 (.A(_00510_),
    .B(net77),
    .Y(n_4235_o_0));
 INVx1_ASAP7_75t_R n_4236 (.A(n_4235_o_0),
    .Y(n_4236_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4237 (.A1(n_4232_o_0),
    .A2(n_4234_o_0),
    .B(net9),
    .C(n_4236_o_0),
    .D(_00948_),
    .Y(n_4237_o_0));
 OAI21xp33_ASAP7_75t_R n_4238 (.A1(n_4227_o_0),
    .A2(n_4228_o_0),
    .B(n_4229_o_0),
    .Y(n_4238_o_0));
 OAI21xp33_ASAP7_75t_R n_4239 (.A1(n_4230_o_0),
    .A2(n_4238_o_0),
    .B(n_4234_o_0),
    .Y(n_4239_o_0));
 AOI211xp5_ASAP7_75t_R n_4240 (.A1(n_4239_o_0),
    .A2(net),
    .B(n_2430_o_0),
    .C(n_4235_o_0),
    .Y(n_4240_o_0));
 NOR2xp67_ASAP7_75t_R n_4241 (.A(n_4237_o_0),
    .B(n_4240_o_0),
    .Y(n_4241_o_0));
 NOR3xp33_ASAP7_75t_R n_4242 (.A(net62),
    .B(net59),
    .C(n_4241_o_0),
    .Y(n_4242_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4243 (.A1(n_4185_o_0),
    .A2(n_4188_o_0),
    .B(n_4189_o_0),
    .C(net77),
    .D(n_4191_o_0),
    .Y(n_4243_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_4244 (.A1(n_4192_o_0),
    .A2(net39),
    .B(n_4198_o_0),
    .C(n_4243_o_0),
    .Y(n_4244_o_0));
 NOR2xp33_ASAP7_75t_R n_4245 (.A(n_4226_o_0),
    .B(n_4241_o_0),
    .Y(n_4245_o_0));
 XNOR2xp5_ASAP7_75t_R n_4246 (.A(_01014_),
    .B(_01019_),
    .Y(n_4246_o_0));
 XNOR2xp5_ASAP7_75t_R n_4247 (.A(_01055_),
    .B(n_4246_o_0),
    .Y(n_4247_o_0));
 XNOR2xp5_ASAP7_75t_R n_4248 (.A(_01054_),
    .B(_01059_),
    .Y(n_4248_o_0));
 XNOR2xp5_ASAP7_75t_R n_4249 (.A(_01063_),
    .B(_01102_),
    .Y(n_4249_o_0));
 XNOR2xp5_ASAP7_75t_R n_4250 (.A(n_4248_o_0),
    .B(n_4249_o_0),
    .Y(n_4250_o_0));
 NOR2xp33_ASAP7_75t_R n_4251 (.A(n_4247_o_0),
    .B(n_4250_o_0),
    .Y(n_4251_o_0));
 AO21x1_ASAP7_75t_R n_4252 (.A1(n_3021_o_0),
    .A2(_00693_),
    .B(_00951_),
    .Y(n_4252_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4253 (.A1(n_4247_o_0),
    .A2(n_4250_o_0),
    .B(n_4251_o_0),
    .C(_00858_),
    .D(n_4252_o_0),
    .Y(n_4253_o_0));
 INVx1_ASAP7_75t_R n_4254 (.A(n_4250_o_0),
    .Y(n_4254_o_0));
 NOR2xp33_ASAP7_75t_R n_4255 (.A(n_4247_o_0),
    .B(n_4254_o_0),
    .Y(n_4255_o_0));
 OAI21xp33_ASAP7_75t_R n_4256 (.A1(_00693_),
    .A2(net39),
    .B(_00951_),
    .Y(n_4256_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4257 (.A1(n_4247_o_0),
    .A2(n_4254_o_0),
    .B(n_4255_o_0),
    .C(net77),
    .D(n_4256_o_0),
    .Y(n_4257_o_0));
 NOR2xp67_ASAP7_75t_R n_4258 (.A(n_4253_o_0),
    .B(n_4257_o_0),
    .Y(n_4258_o_0));
 OAI21xp33_ASAP7_75t_R n_4259 (.A1(n_4244_o_0),
    .A2(n_4245_o_0),
    .B(n_4258_o_0),
    .Y(n_4259_o_0));
 XNOR2xp5_ASAP7_75t_R n_4260 (.A(n_4247_o_0),
    .B(n_4250_o_0),
    .Y(n_4260_o_0));
 INVx1_ASAP7_75t_R n_4261 (.A(n_4260_o_0),
    .Y(n_4261_o_0));
 INVx1_ASAP7_75t_R n_4262 (.A(n_4253_o_0),
    .Y(n_4262_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4263 (.A1(n_4261_o_0),
    .A2(net),
    .B(n_4256_o_0),
    .C(n_4262_o_0),
    .Y(n_4263_o_0));
 OAI21xp33_ASAP7_75t_R n_4264 (.A1(n_4241_o_0),
    .A2(n_4200_o_0),
    .B(n_4263_o_0),
    .Y(n_4264_o_0));
 XNOR2xp5_ASAP7_75t_R n_4265 (.A(_01055_),
    .B(_01059_),
    .Y(n_4265_o_0));
 XNOR2xp5_ASAP7_75t_R n_4266 (.A(_01064_),
    .B(_01103_),
    .Y(n_4266_o_0));
 XNOR2xp5_ASAP7_75t_R n_4267 (.A(n_4265_o_0),
    .B(n_4266_o_0),
    .Y(n_4267_o_0));
 XNOR2xp5_ASAP7_75t_R n_4268 (.A(_01015_),
    .B(_01019_),
    .Y(n_4268_o_0));
 XOR2xp5_ASAP7_75t_R n_4269 (.A(_01056_),
    .B(n_4268_o_0),
    .Y(n_4269_o_0));
 XNOR2xp5_ASAP7_75t_R n_4270 (.A(n_4267_o_0),
    .B(n_4269_o_0),
    .Y(n_4270_o_0));
 NAND2xp33_ASAP7_75t_R n_4271 (.A(_00692_),
    .B(net5),
    .Y(n_4271_o_0));
 OAI21xp33_ASAP7_75t_R n_4272 (.A1(net1),
    .A2(n_4270_o_0),
    .B(n_4271_o_0),
    .Y(n_4272_o_0));
 NAND2xp33_ASAP7_75t_R n_4273 (.A(_00952_),
    .B(n_4272_o_0),
    .Y(n_4273_o_0));
 OA21x2_ASAP7_75t_R n_4274 (.A1(_00952_),
    .A2(n_4272_o_0),
    .B(n_4273_o_0),
    .Y(n_4274_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4275 (.A1(n_4242_o_0),
    .A2(n_4259_o_0),
    .B(n_4264_o_0),
    .C(n_4274_o_0),
    .Y(n_4275_o_0));
 NAND2xp33_ASAP7_75t_R n_4276 (.A(n_2520_o_0),
    .B(n_4272_o_0),
    .Y(n_4276_o_0));
 OAI21xp5_ASAP7_75t_R n_4277 (.A1(n_2520_o_0),
    .A2(n_4272_o_0),
    .B(n_4276_o_0),
    .Y(n_4277_o_0));
 INVx1_ASAP7_75t_R n_4278 (.A(n_4277_o_0),
    .Y(n_4278_o_0));
 NOR2xp67_ASAP7_75t_R n_4279 (.A(n_4244_o_0),
    .B(n_4241_o_0),
    .Y(n_4279_o_0));
 NOR2xp33_ASAP7_75t_R n_4280 (.A(n_4258_o_0),
    .B(n_4279_o_0),
    .Y(n_4280_o_0));
 OAI21xp33_ASAP7_75t_R n_4281 (.A1(net9),
    .A2(n_4217_o_0),
    .B(n_4218_o_0),
    .Y(n_4281_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4282 (.A1(net),
    .A2(n_4217_o_0),
    .B(n_4224_o_0),
    .C(n_4281_o_0),
    .Y(n_4282_o_0));
 NOR2xp33_ASAP7_75t_R n_4283 (.A(n_4241_o_0),
    .B(n_4200_o_0),
    .Y(n_4283_o_0));
 NAND2xp33_ASAP7_75t_R n_4284 (.A(n_4282_o_0),
    .B(n_4283_o_0),
    .Y(n_4284_o_0));
 AOI211xp5_ASAP7_75t_R n_4285 (.A1(n_4227_o_0),
    .A2(n_4228_o_0),
    .B(n_4233_o_0),
    .C(n_4230_o_0),
    .Y(n_4285_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4286 (.A1(n_4230_o_0),
    .A2(n_4238_o_0),
    .B(n_4285_o_0),
    .C(net),
    .D(n_4235_o_0),
    .Y(n_4286_o_0));
 AO21x1_ASAP7_75t_R n_4287 (.A1(_00948_),
    .A2(n_4286_o_0),
    .B(n_4237_o_0),
    .Y(n_4287_o_0));
 OAI21xp33_ASAP7_75t_R n_4288 (.A1(n_4237_o_0),
    .A2(n_4240_o_0),
    .B(n_4226_o_0),
    .Y(n_4288_o_0));
 OAI21xp33_ASAP7_75t_R n_4289 (.A1(n_4226_o_0),
    .A2(n_4287_o_0),
    .B(n_4288_o_0),
    .Y(n_4289_o_0));
 NOR2xp33_ASAP7_75t_R n_4290 (.A(n_4226_o_0),
    .B(n_4287_o_0),
    .Y(n_4290_o_0));
 INVx1_ASAP7_75t_R n_4291 (.A(n_4243_o_0),
    .Y(n_4291_o_0));
 NAND2xp33_ASAP7_75t_R n_4292 (.A(n_4199_o_0),
    .B(n_4291_o_0),
    .Y(n_4292_o_0));
 OAI21xp33_ASAP7_75t_R n_4293 (.A1(n_4290_o_0),
    .A2(n_4292_o_0),
    .B(n_4258_o_0),
    .Y(n_4293_o_0));
 AOI21xp33_ASAP7_75t_R n_4294 (.A1(net62),
    .A2(n_4289_o_0),
    .B(n_4293_o_0),
    .Y(n_4294_o_0));
 AOI21xp33_ASAP7_75t_R n_4295 (.A1(n_4280_o_0),
    .A2(n_4284_o_0),
    .B(n_4294_o_0),
    .Y(n_4295_o_0));
 XNOR2xp5_ASAP7_75t_R n_4296 (.A(_01016_),
    .B(_01056_),
    .Y(n_4296_o_0));
 INVx1_ASAP7_75t_R n_4297 (.A(n_4296_o_0),
    .Y(n_4297_o_0));
 XNOR2xp5_ASAP7_75t_R n_4298 (.A(_01065_),
    .B(_01104_),
    .Y(n_4298_o_0));
 XNOR2xp5_ASAP7_75t_R n_4299 (.A(_01057_),
    .B(n_4298_o_0),
    .Y(n_4299_o_0));
 NOR2xp33_ASAP7_75t_R n_4300 (.A(n_4297_o_0),
    .B(n_4299_o_0),
    .Y(n_4300_o_0));
 NOR2xp33_ASAP7_75t_R n_4301 (.A(_00691_),
    .B(net),
    .Y(n_4301_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4302 (.A1(n_4297_o_0),
    .A2(n_4299_o_0),
    .B(n_4300_o_0),
    .C(net),
    .D(n_4301_o_0),
    .Y(n_4302_o_0));
 NAND2xp33_ASAP7_75t_R n_4303 (.A(_00953_),
    .B(n_4302_o_0),
    .Y(n_4303_o_0));
 OAI21xp5_ASAP7_75t_R n_4304 (.A1(_00953_),
    .A2(n_4302_o_0),
    .B(n_4303_o_0),
    .Y(n_4304_o_0));
 INVx1_ASAP7_75t_R n_4305 (.A(n_4304_o_0),
    .Y(n_4305_o_0));
 OAI21xp33_ASAP7_75t_R n_4306 (.A1(n_4278_o_0),
    .A2(n_4295_o_0),
    .B(n_4305_o_0),
    .Y(n_4306_o_0));
 OAI21xp33_ASAP7_75t_R n_4307 (.A1(_00952_),
    .A2(n_4272_o_0),
    .B(n_4273_o_0),
    .Y(n_4307_o_0));
 OA21x2_ASAP7_75t_R n_4308 (.A1(n_4217_o_0),
    .A2(net2),
    .B(n_4218_o_0),
    .Y(n_4308_o_0));
 AO21x1_ASAP7_75t_R n_4309 (.A1(n_4197_o_0),
    .A2(n_4193_o_0),
    .B(n_2462_o_0),
    .Y(n_4309_o_0));
 XNOR2xp5_ASAP7_75t_R n_4310 (.A(n_4185_o_0),
    .B(n_4196_o_0),
    .Y(n_4310_o_0));
 AOI21xp33_ASAP7_75t_R n_4311 (.A1(n_4192_o_0),
    .A2(net2),
    .B(_00950_),
    .Y(n_4311_o_0));
 OAI21xp33_ASAP7_75t_R n_4312 (.A1(net2),
    .A2(n_4310_o_0),
    .B(n_4311_o_0),
    .Y(n_4312_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4313 (.A1(net2),
    .A2(_00512_),
    .B(n_4309_o_0),
    .C(n_4312_o_0),
    .Y(n_4313_o_0));
 OAI21xp33_ASAP7_75t_R n_4314 (.A1(n_4308_o_0),
    .A2(n_4225_o_0),
    .B(n_4313_o_0),
    .Y(n_4314_o_0));
 NAND2xp33_ASAP7_75t_R n_4315 (.A(n_4287_o_0),
    .B(n_4244_o_0),
    .Y(n_4315_o_0));
 INVx1_ASAP7_75t_R n_4316 (.A(n_4256_o_0),
    .Y(n_4316_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_4317 (.A1(n_3021_o_0),
    .A2(n_4260_o_0),
    .B(n_4316_o_0),
    .C(n_4253_o_0),
    .Y(n_4317_o_0));
 OAI211xp5_ASAP7_75t_R n_4318 (.A1(n_4314_o_0),
    .A2(n_4287_o_0),
    .B(n_4315_o_0),
    .C(n_4317_o_0),
    .Y(n_4318_o_0));
 INVx1_ASAP7_75t_R n_4319 (.A(n_4318_o_0),
    .Y(n_4319_o_0));
 NAND2xp33_ASAP7_75t_R n_4320 (.A(n_4307_o_0),
    .B(n_4319_o_0),
    .Y(n_4320_o_0));
 NOR2xp33_ASAP7_75t_R n_4321 (.A(n_4226_o_0),
    .B(n_4315_o_0),
    .Y(n_4321_o_0));
 NOR2xp67_ASAP7_75t_R n_4322 (.A(n_4282_o_0),
    .B(n_4244_o_0),
    .Y(n_4322_o_0));
 NOR3xp33_ASAP7_75t_R n_4323 (.A(n_4321_o_0),
    .B(n_4322_o_0),
    .C(n_4258_o_0),
    .Y(n_4323_o_0));
 NAND2xp33_ASAP7_75t_R n_4324 (.A(n_4226_o_0),
    .B(n_4287_o_0),
    .Y(n_4324_o_0));
 NOR2xp33_ASAP7_75t_R n_4325 (.A(n_4244_o_0),
    .B(n_4324_o_0),
    .Y(n_4325_o_0));
 INVx1_ASAP7_75t_R n_4326 (.A(n_4325_o_0),
    .Y(n_4326_o_0));
 NAND2xp33_ASAP7_75t_R n_4327 (.A(n_4226_o_0),
    .B(n_4244_o_0),
    .Y(n_4327_o_0));
 AOI211xp5_ASAP7_75t_R n_4328 (.A1(n_4326_o_0),
    .A2(n_4327_o_0),
    .B(n_4274_o_0),
    .C(n_4258_o_0),
    .Y(n_4328_o_0));
 INVx2_ASAP7_75t_R n_4329 (.A(n_4317_o_0),
    .Y(n_4329_o_0));
 NOR2xp33_ASAP7_75t_R n_4330 (.A(n_4244_o_0),
    .B(n_4290_o_0),
    .Y(n_4330_o_0));
 NOR4xp25_ASAP7_75t_R n_4331 (.A(n_4278_o_0),
    .B(n_4329_o_0),
    .C(n_4283_o_0),
    .D(n_4330_o_0),
    .Y(n_4331_o_0));
 AOI211xp5_ASAP7_75t_R n_4332 (.A1(n_4323_o_0),
    .A2(n_4277_o_0),
    .B(n_4328_o_0),
    .C(n_4331_o_0),
    .Y(n_4332_o_0));
 NAND2xp33_ASAP7_75t_R n_4333 (.A(n_4297_o_0),
    .B(n_4299_o_0),
    .Y(n_4333_o_0));
 INVx1_ASAP7_75t_R n_4334 (.A(n_4300_o_0),
    .Y(n_4334_o_0));
 INVx1_ASAP7_75t_R n_4335 (.A(n_4301_o_0),
    .Y(n_4335_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4336 (.A1(n_4333_o_0),
    .A2(n_4334_o_0),
    .B(net2),
    .C(n_4335_o_0),
    .D(n_2386_o_0),
    .Y(n_4336_o_0));
 AOI21xp33_ASAP7_75t_R n_4337 (.A1(n_2386_o_0),
    .A2(n_4302_o_0),
    .B(n_4336_o_0),
    .Y(n_4337_o_0));
 XOR2xp5_ASAP7_75t_R n_4338 (.A(_01017_),
    .B(_01057_),
    .Y(n_4338_o_0));
 XNOR2xp5_ASAP7_75t_R n_4339 (.A(_01058_),
    .B(_01066_),
    .Y(n_4339_o_0));
 XNOR2xp5_ASAP7_75t_R n_4340 (.A(_01105_),
    .B(n_4339_o_0),
    .Y(n_4340_o_0));
 NOR2xp33_ASAP7_75t_R n_4341 (.A(n_4338_o_0),
    .B(n_4340_o_0),
    .Y(n_4341_o_0));
 NOR2xp33_ASAP7_75t_R n_4342 (.A(_00690_),
    .B(net),
    .Y(n_4342_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4343 (.A1(n_4338_o_0),
    .A2(n_4340_o_0),
    .B(n_4341_o_0),
    .C(net),
    .D(n_4342_o_0),
    .Y(n_4343_o_0));
 NAND2xp33_ASAP7_75t_R n_4344 (.A(n_2378_o_0),
    .B(n_4343_o_0),
    .Y(n_4344_o_0));
 OAI21xp33_ASAP7_75t_R n_4345 (.A1(n_4343_o_0),
    .A2(n_2378_o_0),
    .B(n_4344_o_0),
    .Y(n_4345_o_0));
 INVx1_ASAP7_75t_R n_4346 (.A(n_4345_o_0),
    .Y(n_4346_o_0));
 AOI31xp33_ASAP7_75t_R n_4347 (.A1(n_4320_o_0),
    .A2(n_4332_o_0),
    .A3(n_4337_o_0),
    .B(n_4346_o_0),
    .Y(n_4347_o_0));
 OAI21xp33_ASAP7_75t_R n_4348 (.A1(n_4275_o_0),
    .A2(n_4306_o_0),
    .B(n_4347_o_0),
    .Y(n_4348_o_0));
 AOI221xp5_ASAP7_75t_R n_4349 (.A1(_00512_),
    .A2(net2),
    .B1(n_4193_o_0),
    .B2(n_4197_o_0),
    .C(n_2462_o_0),
    .Y(n_4349_o_0));
 NOR2xp33_ASAP7_75t_R n_4350 (.A(n_4282_o_0),
    .B(n_4287_o_0),
    .Y(n_4350_o_0));
 OAI21xp33_ASAP7_75t_R n_4351 (.A1(n_4243_o_0),
    .A2(n_4349_o_0),
    .B(n_4350_o_0),
    .Y(n_4351_o_0));
 NOR2xp33_ASAP7_75t_R n_4352 (.A(n_4313_o_0),
    .B(n_4324_o_0),
    .Y(n_4352_o_0));
 INVx1_ASAP7_75t_R n_4353 (.A(n_4352_o_0),
    .Y(n_4353_o_0));
 OAI211xp5_ASAP7_75t_R n_4354 (.A1(n_4308_o_0),
    .A2(n_4225_o_0),
    .B(n_4241_o_0),
    .C(n_4244_o_0),
    .Y(n_4354_o_0));
 INVx1_ASAP7_75t_R n_4355 (.A(n_4354_o_0),
    .Y(n_4355_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4356 (.A1(n_4239_o_0),
    .A2(net),
    .B(n_4235_o_0),
    .C(n_2430_o_0),
    .Y(n_4356_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4357 (.A1(n_4230_o_0),
    .A2(n_4238_o_0),
    .B(n_4285_o_0),
    .C(net),
    .Y(n_4357_o_0));
 OAI211xp5_ASAP7_75t_R n_4358 (.A1(_00510_),
    .A2(net),
    .B(n_4357_o_0),
    .C(_00948_),
    .Y(n_4358_o_0));
 INVx1_ASAP7_75t_R n_4359 (.A(n_4225_o_0),
    .Y(n_4359_o_0));
 AOI33xp33_ASAP7_75t_R n_4360 (.A1(n_4356_o_0),
    .A2(n_4282_o_0),
    .A3(n_4358_o_0),
    .B1(n_4287_o_0),
    .B2(n_4359_o_0),
    .B3(n_4281_o_0),
    .Y(n_4360_o_0));
 OAI21xp33_ASAP7_75t_R n_4361 (.A1(n_4244_o_0),
    .A2(n_4360_o_0),
    .B(n_4263_o_0),
    .Y(n_4361_o_0));
 NOR2xp33_ASAP7_75t_R n_4362 (.A(n_4355_o_0),
    .B(n_4361_o_0),
    .Y(n_4362_o_0));
 AOI31xp33_ASAP7_75t_R n_4363 (.A1(n_4351_o_0),
    .A2(n_4353_o_0),
    .A3(net27),
    .B(n_4362_o_0),
    .Y(n_4363_o_0));
 NAND2xp33_ASAP7_75t_R n_4364 (.A(n_4244_o_0),
    .B(n_4241_o_0),
    .Y(n_4364_o_0));
 INVx1_ASAP7_75t_R n_4365 (.A(n_4364_o_0),
    .Y(n_4365_o_0));
 NOR2xp33_ASAP7_75t_R n_4366 (.A(n_4226_o_0),
    .B(n_4241_o_0),
    .Y(n_4366_o_0));
 NAND2xp33_ASAP7_75t_R n_4367 (.A(n_4241_o_0),
    .B(n_4200_o_0),
    .Y(n_4367_o_0));
 NAND2xp33_ASAP7_75t_R n_4368 (.A(n_4226_o_0),
    .B(n_4287_o_0),
    .Y(n_4368_o_0));
 NAND3xp33_ASAP7_75t_R n_4369 (.A(n_4367_o_0),
    .B(n_4368_o_0),
    .C(n_4263_o_0),
    .Y(n_4369_o_0));
 OAI31xp33_ASAP7_75t_R n_4370 (.A1(n_4365_o_0),
    .A2(n_4366_o_0),
    .A3(n_4329_o_0),
    .B(n_4369_o_0),
    .Y(n_4370_o_0));
 INVx1_ASAP7_75t_R n_4371 (.A(n_4370_o_0),
    .Y(n_4371_o_0));
 OAI22xp33_ASAP7_75t_R n_4372 (.A1(n_4363_o_0),
    .A2(n_4274_o_0),
    .B1(n_4278_o_0),
    .B2(n_4371_o_0),
    .Y(n_4372_o_0));
 NAND4xp25_ASAP7_75t_R n_4373 (.A(n_4221_o_0),
    .B(n_4207_o_0),
    .C(n_4222_o_0),
    .D(n_4203_o_0),
    .Y(n_4373_o_0));
 AOI211xp5_ASAP7_75t_R n_4374 (.A1(n_4373_o_0),
    .A2(n_4216_o_0),
    .B(net2),
    .C(n_2445_o_0),
    .Y(n_4374_o_0));
 NOR3xp33_ASAP7_75t_R n_4375 (.A(n_2445_o_0),
    .B(net),
    .C(_00509_),
    .Y(n_4375_o_0));
 OAI311xp33_ASAP7_75t_R n_4376 (.A1(n_4225_o_0),
    .A2(n_4374_o_0),
    .A3(n_4375_o_0),
    .B1(n_4358_o_0),
    .C1(n_4356_o_0),
    .Y(n_4376_o_0));
 OAI211xp5_ASAP7_75t_R n_4377 (.A1(n_4243_o_0),
    .A2(n_4349_o_0),
    .B(n_4288_o_0),
    .C(n_4376_o_0),
    .Y(n_4377_o_0));
 NAND2xp33_ASAP7_75t_R n_4378 (.A(n_4263_o_0),
    .B(n_4377_o_0),
    .Y(n_4378_o_0));
 NOR2xp33_ASAP7_75t_R n_4379 (.A(n_4226_o_0),
    .B(n_4200_o_0),
    .Y(n_4379_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4380 (.A1(n_4288_o_0),
    .A2(n_4376_o_0),
    .B(n_4313_o_0),
    .C(n_4317_o_0),
    .Y(n_4380_o_0));
 OAI211xp5_ASAP7_75t_R n_4381 (.A1(n_4378_o_0),
    .A2(n_4379_o_0),
    .B(n_4380_o_0),
    .C(n_4274_o_0),
    .Y(n_4381_o_0));
 AOI22xp33_ASAP7_75t_R n_4382 (.A1(n_4291_o_0),
    .A2(n_4199_o_0),
    .B1(n_4287_o_0),
    .B2(n_4226_o_0),
    .Y(n_4382_o_0));
 INVx1_ASAP7_75t_R n_4383 (.A(n_4382_o_0),
    .Y(n_4383_o_0));
 NOR2xp33_ASAP7_75t_R n_4384 (.A(n_4317_o_0),
    .B(n_4383_o_0),
    .Y(n_4384_o_0));
 AOI21xp33_ASAP7_75t_R n_4385 (.A1(n_4200_o_0),
    .A2(n_4289_o_0),
    .B(n_4329_o_0),
    .Y(n_4385_o_0));
 OAI21xp33_ASAP7_75t_R n_4386 (.A1(n_4324_o_0),
    .A2(n_4313_o_0),
    .B(n_4385_o_0),
    .Y(n_4386_o_0));
 OAI31xp33_ASAP7_75t_R n_4387 (.A1(n_4258_o_0),
    .A2(n_4350_o_0),
    .A3(net62),
    .B(n_4386_o_0),
    .Y(n_4387_o_0));
 OAI21xp33_ASAP7_75t_R n_4388 (.A1(n_4384_o_0),
    .A2(n_4387_o_0),
    .B(n_4307_o_0),
    .Y(n_4388_o_0));
 NAND2xp33_ASAP7_75t_R n_4389 (.A(_00954_),
    .B(n_4343_o_0),
    .Y(n_4389_o_0));
 OAI21xp33_ASAP7_75t_R n_4390 (.A1(_00954_),
    .A2(n_4343_o_0),
    .B(n_4389_o_0),
    .Y(n_4390_o_0));
 INVx1_ASAP7_75t_R n_4391 (.A(n_4390_o_0),
    .Y(n_4391_o_0));
 AOI31xp33_ASAP7_75t_R n_4392 (.A1(n_4381_o_0),
    .A2(n_4388_o_0),
    .A3(n_4337_o_0),
    .B(n_4391_o_0),
    .Y(n_4392_o_0));
 OAI21xp33_ASAP7_75t_R n_4393 (.A1(n_4304_o_0),
    .A2(n_4372_o_0),
    .B(n_4392_o_0),
    .Y(n_4393_o_0));
 XOR2xp5_ASAP7_75t_R n_4394 (.A(_01018_),
    .B(_01058_),
    .Y(n_4394_o_0));
 XNOR2xp5_ASAP7_75t_R n_4395 (.A(_01059_),
    .B(_01067_),
    .Y(n_4395_o_0));
 XNOR2xp5_ASAP7_75t_R n_4396 (.A(_01106_),
    .B(n_4395_o_0),
    .Y(n_4396_o_0));
 NOR2xp33_ASAP7_75t_R n_4397 (.A(n_4394_o_0),
    .B(n_4396_o_0),
    .Y(n_4397_o_0));
 NOR2xp33_ASAP7_75t_R n_4398 (.A(_00689_),
    .B(net),
    .Y(n_4398_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4399 (.A1(n_4394_o_0),
    .A2(n_4396_o_0),
    .B(n_4397_o_0),
    .C(net),
    .D(n_4398_o_0),
    .Y(n_4399_o_0));
 NAND2xp33_ASAP7_75t_R n_4400 (.A(_00955_),
    .B(n_4399_o_0),
    .Y(n_4400_o_0));
 OAI21xp33_ASAP7_75t_R n_4401 (.A1(_00955_),
    .A2(n_4399_o_0),
    .B(n_4400_o_0),
    .Y(n_4401_o_0));
 INVx1_ASAP7_75t_R n_4402 (.A(n_4401_o_0),
    .Y(n_4402_o_0));
 OAI21xp33_ASAP7_75t_R n_4403 (.A1(n_4287_o_0),
    .A2(n_4282_o_0),
    .B(n_4244_o_0),
    .Y(n_4403_o_0));
 NAND2xp33_ASAP7_75t_R n_4404 (.A(n_4317_o_0),
    .B(n_4403_o_0),
    .Y(n_4404_o_0));
 AOI221xp5_ASAP7_75t_R n_4405 (.A1(_00512_),
    .A2(net2),
    .B1(n_4193_o_0),
    .B2(n_4197_o_0),
    .C(n_2462_o_0),
    .Y(n_4405_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4406 (.A1(n_4310_o_0),
    .A2(net2),
    .B(n_4311_o_0),
    .C(n_4405_o_0),
    .Y(n_4406_o_0));
 AOI211xp5_ASAP7_75t_R n_4407 (.A1(n_4281_o_0),
    .A2(n_4359_o_0),
    .B(n_4241_o_0),
    .C(n_4406_o_0),
    .Y(n_4407_o_0));
 INVx1_ASAP7_75t_R n_4408 (.A(n_4324_o_0),
    .Y(n_4408_o_0));
 NAND3xp33_ASAP7_75t_R n_4409 (.A(n_4408_o_0),
    .B(n_4329_o_0),
    .C(n_4200_o_0),
    .Y(n_4409_o_0));
 OAI211xp5_ASAP7_75t_R n_4410 (.A1(n_4404_o_0),
    .A2(n_4407_o_0),
    .B(n_4409_o_0),
    .C(n_4307_o_0),
    .Y(n_4410_o_0));
 INVx1_ASAP7_75t_R n_4411 (.A(n_4350_o_0),
    .Y(n_4411_o_0));
 OAI21xp33_ASAP7_75t_R n_4412 (.A1(n_4313_o_0),
    .A2(n_4411_o_0),
    .B(n_4263_o_0),
    .Y(n_4412_o_0));
 AOI21xp33_ASAP7_75t_R n_4413 (.A1(n_4317_o_0),
    .A2(n_4325_o_0),
    .B(n_4307_o_0),
    .Y(n_4413_o_0));
 OAI21xp33_ASAP7_75t_R n_4414 (.A1(n_4407_o_0),
    .A2(n_4412_o_0),
    .B(n_4413_o_0),
    .Y(n_4414_o_0));
 NAND3xp33_ASAP7_75t_R n_4415 (.A(n_4410_o_0),
    .B(n_4414_o_0),
    .C(n_4305_o_0),
    .Y(n_4415_o_0));
 OAI21xp33_ASAP7_75t_R n_4416 (.A1(n_4241_o_0),
    .A2(net47),
    .B(n_4329_o_0),
    .Y(n_4416_o_0));
 AOI21xp33_ASAP7_75t_R n_4417 (.A1(net47),
    .A2(n_4324_o_0),
    .B(n_4416_o_0),
    .Y(n_4417_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4418 (.A1(n_4383_o_0),
    .A2(n_4364_o_0),
    .B(n_4263_o_0),
    .C(n_4307_o_0),
    .Y(n_4418_o_0));
 NOR2xp33_ASAP7_75t_R n_4419 (.A(n_4292_o_0),
    .B(n_4245_o_0),
    .Y(n_4419_o_0));
 AOI21xp33_ASAP7_75t_R n_4420 (.A1(n_4281_o_0),
    .A2(n_4359_o_0),
    .B(n_4406_o_0),
    .Y(n_4420_o_0));
 NOR3xp33_ASAP7_75t_R n_4421 (.A(n_4419_o_0),
    .B(n_4420_o_0),
    .C(net27),
    .Y(n_4421_o_0));
 AOI21xp33_ASAP7_75t_R n_4422 (.A1(n_4244_o_0),
    .A2(n_4360_o_0),
    .B(n_4258_o_0),
    .Y(n_4422_o_0));
 NOR2xp33_ASAP7_75t_R n_4423 (.A(net59),
    .B(net47),
    .Y(n_4423_o_0));
 OAI21xp33_ASAP7_75t_R n_4424 (.A1(n_4329_o_0),
    .A2(n_4423_o_0),
    .B(n_4337_o_0),
    .Y(n_4424_o_0));
 NAND2xp33_ASAP7_75t_R n_4425 (.A(n_4304_o_0),
    .B(n_4307_o_0),
    .Y(n_4425_o_0));
 OAI21xp33_ASAP7_75t_R n_4426 (.A1(n_4422_o_0),
    .A2(n_4424_o_0),
    .B(n_4425_o_0),
    .Y(n_4426_o_0));
 OAI31xp33_ASAP7_75t_R n_4427 (.A1(n_4417_o_0),
    .A2(n_4418_o_0),
    .A3(n_4421_o_0),
    .B(n_4426_o_0),
    .Y(n_4427_o_0));
 AOI21xp33_ASAP7_75t_R n_4428 (.A1(n_4415_o_0),
    .A2(n_4427_o_0),
    .B(n_4345_o_0),
    .Y(n_4428_o_0));
 OAI21xp33_ASAP7_75t_R n_4429 (.A1(n_4244_o_0),
    .A2(n_4360_o_0),
    .B(n_4317_o_0),
    .Y(n_4429_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4430 (.A1(n_4351_o_0),
    .A2(net27),
    .B(n_4429_o_0),
    .C(n_4278_o_0),
    .Y(n_4430_o_0));
 NAND2xp33_ASAP7_75t_R n_4431 (.A(n_4282_o_0),
    .B(n_4287_o_0),
    .Y(n_4431_o_0));
 NOR3xp33_ASAP7_75t_R n_4432 (.A(n_4431_o_0),
    .B(n_4313_o_0),
    .C(n_4317_o_0),
    .Y(n_4432_o_0));
 AOI211xp5_ASAP7_75t_R n_4433 (.A1(n_4319_o_0),
    .A2(n_4307_o_0),
    .B(n_4430_o_0),
    .C(n_4432_o_0),
    .Y(n_4433_o_0));
 NOR2xp33_ASAP7_75t_R n_4434 (.A(n_4313_o_0),
    .B(n_4411_o_0),
    .Y(n_4434_o_0));
 NAND2xp33_ASAP7_75t_R n_4435 (.A(n_4282_o_0),
    .B(n_4200_o_0),
    .Y(n_4435_o_0));
 NAND2xp33_ASAP7_75t_R n_4436 (.A(n_4435_o_0),
    .B(n_4422_o_0),
    .Y(n_4436_o_0));
 OAI31xp33_ASAP7_75t_R n_4437 (.A1(n_4434_o_0),
    .A2(n_4279_o_0),
    .A3(n_4329_o_0),
    .B(n_4436_o_0),
    .Y(n_4437_o_0));
 AOI21xp33_ASAP7_75t_R n_4438 (.A1(n_4226_o_0),
    .A2(n_4287_o_0),
    .B(n_4313_o_0),
    .Y(n_4438_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4439 (.A1(n_4408_o_0),
    .A2(n_4200_o_0),
    .B(n_4438_o_0),
    .C(n_4329_o_0),
    .Y(n_4439_o_0));
 AOI21xp33_ASAP7_75t_R n_4440 (.A1(n_4259_o_0),
    .A2(n_4439_o_0),
    .B(n_4307_o_0),
    .Y(n_4440_o_0));
 AOI211xp5_ASAP7_75t_R n_4441 (.A1(n_4437_o_0),
    .A2(n_4307_o_0),
    .B(n_4337_o_0),
    .C(n_4440_o_0),
    .Y(n_4441_o_0));
 AOI211xp5_ASAP7_75t_R n_4442 (.A1(n_4433_o_0),
    .A2(n_4304_o_0),
    .B(n_4441_o_0),
    .C(n_4390_o_0),
    .Y(n_4442_o_0));
 OAI21xp33_ASAP7_75t_R n_4443 (.A1(n_4428_o_0),
    .A2(n_4442_o_0),
    .B(n_4402_o_0),
    .Y(n_4443_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4444 (.A1(n_4348_o_0),
    .A2(n_4393_o_0),
    .B(n_4402_o_0),
    .C(n_4443_o_0),
    .Y(n_4444_o_0));
 AOI21xp33_ASAP7_75t_R n_4445 (.A1(n_4244_o_0),
    .A2(n_4226_o_0),
    .B(n_4329_o_0),
    .Y(n_4445_o_0));
 OAI21xp33_ASAP7_75t_R n_4446 (.A1(net47),
    .A2(n_4245_o_0),
    .B(n_4445_o_0),
    .Y(n_4446_o_0));
 NOR2xp33_ASAP7_75t_R n_4447 (.A(n_4287_o_0),
    .B(n_4244_o_0),
    .Y(n_4447_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4448 (.A1(n_4258_o_0),
    .A2(n_4379_o_0),
    .B(n_4446_o_0),
    .C(n_4447_o_0),
    .Y(n_4448_o_0));
 INVx1_ASAP7_75t_R n_4449 (.A(n_4448_o_0),
    .Y(n_4449_o_0));
 NOR3xp33_ASAP7_75t_R n_4450 (.A(n_4200_o_0),
    .B(n_4257_o_0),
    .C(n_4253_o_0),
    .Y(n_4450_o_0));
 INVx1_ASAP7_75t_R n_4451 (.A(n_4366_o_0),
    .Y(n_4451_o_0));
 AOI21xp33_ASAP7_75t_R n_4452 (.A1(n_4450_o_0),
    .A2(n_4451_o_0),
    .B(n_4304_o_0),
    .Y(n_4452_o_0));
 NOR2xp33_ASAP7_75t_R n_4453 (.A(n_4226_o_0),
    .B(n_4287_o_0),
    .Y(n_4453_o_0));
 INVx1_ASAP7_75t_R n_4454 (.A(n_4453_o_0),
    .Y(n_4454_o_0));
 NOR3xp33_ASAP7_75t_R n_4455 (.A(n_4352_o_0),
    .B(n_4279_o_0),
    .C(n_4258_o_0),
    .Y(n_4455_o_0));
 AOI31xp33_ASAP7_75t_R n_4456 (.A1(net62),
    .A2(n_4454_o_0),
    .A3(net27),
    .B(n_4455_o_0),
    .Y(n_4456_o_0));
 AOI22xp33_ASAP7_75t_R n_4457 (.A1(n_4449_o_0),
    .A2(n_4337_o_0),
    .B1(n_4452_o_0),
    .B2(n_4456_o_0),
    .Y(n_4457_o_0));
 AOI211xp5_ASAP7_75t_R n_4458 (.A1(n_4358_o_0),
    .A2(n_4356_o_0),
    .B(n_4308_o_0),
    .C(n_4225_o_0),
    .Y(n_4458_o_0));
 AOI211xp5_ASAP7_75t_R n_4459 (.A1(n_4359_o_0),
    .A2(n_4281_o_0),
    .B(n_4240_o_0),
    .C(n_4237_o_0),
    .Y(n_4459_o_0));
 AOI211xp5_ASAP7_75t_R n_4460 (.A1(n_4291_o_0),
    .A2(n_4199_o_0),
    .B(n_4458_o_0),
    .C(n_4459_o_0),
    .Y(n_4460_o_0));
 NOR3xp33_ASAP7_75t_R n_4461 (.A(n_4355_o_0),
    .B(n_4329_o_0),
    .C(n_4460_o_0),
    .Y(n_4461_o_0));
 INVx1_ASAP7_75t_R n_4462 (.A(n_4438_o_0),
    .Y(n_4462_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4463 (.A1(n_4226_o_0),
    .A2(n_4287_o_0),
    .B(n_4200_o_0),
    .C(n_4317_o_0),
    .Y(n_4463_o_0));
 AO21x1_ASAP7_75t_R n_4464 (.A1(n_2386_o_0),
    .A2(n_4302_o_0),
    .B(n_4336_o_0),
    .Y(n_4464_o_0));
 AO21x1_ASAP7_75t_R n_4465 (.A1(n_4462_o_0),
    .A2(n_4463_o_0),
    .B(n_4464_o_0),
    .Y(n_4465_o_0));
 OAI21xp33_ASAP7_75t_R n_4466 (.A1(n_4461_o_0),
    .A2(n_4465_o_0),
    .B(n_4345_o_0),
    .Y(n_4466_o_0));
 NAND2xp33_ASAP7_75t_R n_4467 (.A(net47),
    .B(n_4258_o_0),
    .Y(n_4467_o_0));
 OAI221xp5_ASAP7_75t_R n_4468 (.A1(n_4383_o_0),
    .A2(n_4263_o_0),
    .B1(n_4289_o_0),
    .B2(n_4467_o_0),
    .C(n_4409_o_0),
    .Y(n_4468_o_0));
 AOI311xp33_ASAP7_75t_R n_4469 (.A1(n_4241_o_0),
    .A2(net47),
    .A3(n_4329_o_0),
    .B(n_4337_o_0),
    .C(n_4468_o_0),
    .Y(n_4469_o_0));
 XNOR2xp5_ASAP7_75t_R n_4470 (.A(_00955_),
    .B(n_4399_o_0),
    .Y(n_4470_o_0));
 OAI21xp33_ASAP7_75t_R n_4471 (.A1(n_4466_o_0),
    .A2(n_4469_o_0),
    .B(n_4470_o_0),
    .Y(n_4471_o_0));
 AOI21xp33_ASAP7_75t_R n_4472 (.A1(n_4390_o_0),
    .A2(n_4457_o_0),
    .B(n_4471_o_0),
    .Y(n_4472_o_0));
 OAI21xp33_ASAP7_75t_R n_4473 (.A1(net59),
    .A2(n_4200_o_0),
    .B(n_4317_o_0),
    .Y(n_4473_o_0));
 INVx1_ASAP7_75t_R n_4474 (.A(n_4421_o_0),
    .Y(n_4474_o_0));
 AOI21xp33_ASAP7_75t_R n_4475 (.A1(n_4287_o_0),
    .A2(n_4282_o_0),
    .B(n_4244_o_0),
    .Y(n_4475_o_0));
 OAI31xp33_ASAP7_75t_R n_4476 (.A1(n_4475_o_0),
    .A2(n_4365_o_0),
    .A3(n_4258_o_0),
    .B(n_4305_o_0),
    .Y(n_4476_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4477 (.A1(n_4315_o_0),
    .A2(n_4385_o_0),
    .B(n_4476_o_0),
    .C(n_4390_o_0),
    .Y(n_4477_o_0));
 AOI31xp33_ASAP7_75t_R n_4478 (.A1(n_4473_o_0),
    .A2(n_4474_o_0),
    .A3(n_4304_o_0),
    .B(n_4477_o_0),
    .Y(n_4478_o_0));
 OAI21xp33_ASAP7_75t_R n_4479 (.A1(n_4313_o_0),
    .A2(n_4431_o_0),
    .B(n_4385_o_0),
    .Y(n_4479_o_0));
 OAI31xp33_ASAP7_75t_R n_4480 (.A1(n_4365_o_0),
    .A2(n_4382_o_0),
    .A3(n_4258_o_0),
    .B(n_4479_o_0),
    .Y(n_4480_o_0));
 AOI21xp33_ASAP7_75t_R n_4481 (.A1(n_4282_o_0),
    .A2(n_4241_o_0),
    .B(n_4244_o_0),
    .Y(n_4481_o_0));
 AOI21xp33_ASAP7_75t_R n_4482 (.A1(n_4329_o_0),
    .A2(n_4481_o_0),
    .B(n_4337_o_0),
    .Y(n_4482_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4483 (.A1(net62),
    .A2(net59),
    .B(n_4293_o_0),
    .C(n_4482_o_0),
    .Y(n_4483_o_0));
 INVx1_ASAP7_75t_R n_4484 (.A(n_4483_o_0),
    .Y(n_4484_o_0));
 AOI211xp5_ASAP7_75t_R n_4485 (.A1(n_4480_o_0),
    .A2(n_4304_o_0),
    .B(n_4390_o_0),
    .C(n_4484_o_0),
    .Y(n_4485_o_0));
 NOR3xp33_ASAP7_75t_R n_4486 (.A(n_4478_o_0),
    .B(n_4485_o_0),
    .C(n_4401_o_0),
    .Y(n_4486_o_0));
 NOR2xp33_ASAP7_75t_R n_4487 (.A(n_4317_o_0),
    .B(n_4420_o_0),
    .Y(n_4487_o_0));
 NAND2xp33_ASAP7_75t_R n_4488 (.A(n_4368_o_0),
    .B(n_4487_o_0),
    .Y(n_4488_o_0));
 NOR3xp33_ASAP7_75t_R n_4489 (.A(n_4258_o_0),
    .B(net82),
    .C(net47),
    .Y(n_4489_o_0));
 OAI221xp5_ASAP7_75t_R n_4490 (.A1(n_4241_o_0),
    .A2(net47),
    .B1(n_4292_o_0),
    .B2(n_4245_o_0),
    .C(n_4329_o_0),
    .Y(n_4490_o_0));
 INVx1_ASAP7_75t_R n_4491 (.A(n_4490_o_0),
    .Y(n_4491_o_0));
 OAI21xp33_ASAP7_75t_R n_4492 (.A1(n_4380_o_0),
    .A2(n_4330_o_0),
    .B(n_4337_o_0),
    .Y(n_4492_o_0));
 OAI31xp33_ASAP7_75t_R n_4493 (.A1(n_4489_o_0),
    .A2(n_4491_o_0),
    .A3(n_4492_o_0),
    .B(n_4390_o_0),
    .Y(n_4493_o_0));
 OAI31xp33_ASAP7_75t_R n_4494 (.A1(net47),
    .A2(n_4431_o_0),
    .A3(net27),
    .B(n_4305_o_0),
    .Y(n_4494_o_0));
 INVx1_ASAP7_75t_R n_4495 (.A(n_4422_o_0),
    .Y(n_4495_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4496 (.A1(n_4453_o_0),
    .A2(n_4279_o_0),
    .B(n_4317_o_0),
    .C(n_4464_o_0),
    .Y(n_4496_o_0));
 OAI21xp33_ASAP7_75t_R n_4497 (.A1(n_4279_o_0),
    .A2(n_4495_o_0),
    .B(n_4496_o_0),
    .Y(n_4497_o_0));
 OAI211xp5_ASAP7_75t_R n_4498 (.A1(n_4494_o_0),
    .A2(n_4461_o_0),
    .B(n_4497_o_0),
    .C(n_4345_o_0),
    .Y(n_4498_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4499 (.A1(n_4452_o_0),
    .A2(n_4488_o_0),
    .B(n_4493_o_0),
    .C(n_4498_o_0),
    .Y(n_4499_o_0));
 NOR2xp33_ASAP7_75t_R n_4500 (.A(net82),
    .B(net62),
    .Y(n_4500_o_0));
 NAND2xp33_ASAP7_75t_R n_4501 (.A(n_4241_o_0),
    .B(n_4420_o_0),
    .Y(n_4501_o_0));
 OAI211xp5_ASAP7_75t_R n_4502 (.A1(n_4313_o_0),
    .A2(n_4411_o_0),
    .B(n_4501_o_0),
    .C(n_4263_o_0),
    .Y(n_4502_o_0));
 OAI31xp33_ASAP7_75t_R n_4503 (.A1(n_4305_o_0),
    .A2(n_4500_o_0),
    .A3(n_4329_o_0),
    .B(n_4502_o_0),
    .Y(n_4503_o_0));
 INVx1_ASAP7_75t_R n_4504 (.A(n_4470_o_0),
    .Y(n_4504_o_0));
 AOI21xp33_ASAP7_75t_R n_4505 (.A1(n_4390_o_0),
    .A2(n_4503_o_0),
    .B(n_4504_o_0),
    .Y(n_4505_o_0));
 INVx1_ASAP7_75t_R n_4506 (.A(n_4501_o_0),
    .Y(n_4506_o_0));
 OAI211xp5_ASAP7_75t_R n_4507 (.A1(n_4506_o_0),
    .A2(n_4264_o_0),
    .B(n_4429_o_0),
    .C(n_4337_o_0),
    .Y(n_4507_o_0));
 NAND2xp33_ASAP7_75t_R n_4508 (.A(n_4263_o_0),
    .B(n_4367_o_0),
    .Y(n_4508_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4509 (.A1(net47),
    .A2(n_4245_o_0),
    .B(n_4445_o_0),
    .C(n_4304_o_0),
    .Y(n_4509_o_0));
 OAI21xp33_ASAP7_75t_R n_4510 (.A1(n_4508_o_0),
    .A2(n_4352_o_0),
    .B(n_4509_o_0),
    .Y(n_4510_o_0));
 NAND3xp33_ASAP7_75t_R n_4511 (.A(n_4507_o_0),
    .B(n_4510_o_0),
    .C(n_4345_o_0),
    .Y(n_4511_o_0));
 AOI21xp33_ASAP7_75t_R n_4512 (.A1(n_4505_o_0),
    .A2(n_4511_o_0),
    .B(n_4274_o_0),
    .Y(n_4512_o_0));
 OAI21xp33_ASAP7_75t_R n_4513 (.A1(n_4401_o_0),
    .A2(n_4499_o_0),
    .B(n_4512_o_0),
    .Y(n_4513_o_0));
 OAI31xp33_ASAP7_75t_R n_4514 (.A1(n_4278_o_0),
    .A2(n_4472_o_0),
    .A3(n_4486_o_0),
    .B(n_4513_o_0),
    .Y(n_4514_o_0));
 INVx1_ASAP7_75t_R n_4515 (.A(n_4445_o_0),
    .Y(n_4515_o_0));
 INVx1_ASAP7_75t_R n_4516 (.A(n_4351_o_0),
    .Y(n_4516_o_0));
 OAI31xp33_ASAP7_75t_R n_4517 (.A1(n_4287_o_0),
    .A2(net59),
    .A3(n_4200_o_0),
    .B(n_4263_o_0),
    .Y(n_4517_o_0));
 OA21x2_ASAP7_75t_R n_4518 (.A1(n_4517_o_0),
    .A2(n_4447_o_0),
    .B(n_4274_o_0),
    .Y(n_4518_o_0));
 OAI21xp33_ASAP7_75t_R n_4519 (.A1(n_4515_o_0),
    .A2(n_4516_o_0),
    .B(n_4518_o_0),
    .Y(n_4519_o_0));
 OAI21xp33_ASAP7_75t_R n_4520 (.A1(net62),
    .A2(n_4289_o_0),
    .B(n_4385_o_0),
    .Y(n_4520_o_0));
 OAI211xp5_ASAP7_75t_R n_4521 (.A1(net59),
    .A2(n_4200_o_0),
    .B(n_4329_o_0),
    .C(n_4241_o_0),
    .Y(n_4521_o_0));
 AO21x1_ASAP7_75t_R n_4522 (.A1(n_4520_o_0),
    .A2(n_4521_o_0),
    .B(n_4277_o_0),
    .Y(n_4522_o_0));
 OAI211xp5_ASAP7_75t_R n_4523 (.A1(n_4313_o_0),
    .A2(n_4431_o_0),
    .B(n_4367_o_0),
    .C(n_4317_o_0),
    .Y(n_4523_o_0));
 AOI21xp33_ASAP7_75t_R n_4524 (.A1(net82),
    .A2(n_4258_o_0),
    .B(net47),
    .Y(n_4524_o_0));
 OAI31xp33_ASAP7_75t_R n_4525 (.A1(n_4524_o_0),
    .A2(n_4419_o_0),
    .A3(n_4277_o_0),
    .B(n_4304_o_0),
    .Y(n_4525_o_0));
 AOI321xp33_ASAP7_75t_R n_4526 (.A1(n_4523_o_0),
    .A2(n_4517_o_0),
    .A3(n_4274_o_0),
    .B1(n_4516_o_0),
    .B2(n_4329_o_0),
    .C(n_4525_o_0),
    .Y(n_4526_o_0));
 AOI31xp33_ASAP7_75t_R n_4527 (.A1(n_4464_o_0),
    .A2(n_4519_o_0),
    .A3(n_4522_o_0),
    .B(n_4526_o_0),
    .Y(n_4527_o_0));
 OAI21xp33_ASAP7_75t_R n_4528 (.A1(n_4402_o_0),
    .A2(n_4527_o_0),
    .B(n_4391_o_0),
    .Y(n_4528_o_0));
 AOI31xp33_ASAP7_75t_R n_4529 (.A1(n_4258_o_0),
    .A2(n_4314_o_0),
    .A3(n_4368_o_0),
    .B(n_4277_o_0),
    .Y(n_4529_o_0));
 NAND2xp33_ASAP7_75t_R n_4530 (.A(n_4406_o_0),
    .B(n_4289_o_0),
    .Y(n_4530_o_0));
 AOI21xp33_ASAP7_75t_R n_4531 (.A1(n_4351_o_0),
    .A2(n_4530_o_0),
    .B(n_4263_o_0),
    .Y(n_4531_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4532 (.A1(n_4462_o_0),
    .A2(n_4487_o_0),
    .B(n_4531_o_0),
    .C(n_4274_o_0),
    .Y(n_4532_o_0));
 NAND2xp33_ASAP7_75t_R n_4533 (.A(n_4304_o_0),
    .B(n_4532_o_0),
    .Y(n_4533_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4534 (.A1(net47),
    .A2(net59),
    .B(n_4258_o_0),
    .C(n_4529_o_0),
    .D(n_4533_o_0),
    .Y(n_4534_o_0));
 AOI21xp33_ASAP7_75t_R n_4535 (.A1(n_4435_o_0),
    .A2(n_4422_o_0),
    .B(n_4307_o_0),
    .Y(n_4535_o_0));
 AOI21xp33_ASAP7_75t_R n_4536 (.A1(n_4244_o_0),
    .A2(net59),
    .B(n_4279_o_0),
    .Y(n_4536_o_0));
 NAND2xp33_ASAP7_75t_R n_4537 (.A(net27),
    .B(n_4536_o_0),
    .Y(n_4537_o_0));
 OAI21xp33_ASAP7_75t_R n_4538 (.A1(n_4380_o_0),
    .A2(n_4407_o_0),
    .B(n_4278_o_0),
    .Y(n_4538_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4539 (.A1(n_4263_o_0),
    .A2(n_4423_o_0),
    .B(n_4538_o_0),
    .C(n_4464_o_0),
    .Y(n_4539_o_0));
 AOI21xp33_ASAP7_75t_R n_4540 (.A1(n_4535_o_0),
    .A2(n_4537_o_0),
    .B(n_4539_o_0),
    .Y(n_4540_o_0));
 NOR3xp33_ASAP7_75t_R n_4541 (.A(n_4534_o_0),
    .B(n_4540_o_0),
    .C(n_4401_o_0),
    .Y(n_4541_o_0));
 AOI21xp33_ASAP7_75t_R n_4542 (.A1(net62),
    .A2(net82),
    .B(n_4495_o_0),
    .Y(n_4542_o_0));
 OAI21xp33_ASAP7_75t_R n_4543 (.A1(n_4322_o_0),
    .A2(n_4523_o_0),
    .B(n_4278_o_0),
    .Y(n_4543_o_0));
 NOR2xp33_ASAP7_75t_R n_4544 (.A(n_2520_o_0),
    .B(n_4272_o_0),
    .Y(n_4544_o_0));
 OAI21xp33_ASAP7_75t_R n_4545 (.A1(n_4287_o_0),
    .A2(n_4226_o_0),
    .B(n_4244_o_0),
    .Y(n_4545_o_0));
 INVx1_ASAP7_75t_R n_4546 (.A(n_4545_o_0),
    .Y(n_4546_o_0));
 OAI211xp5_ASAP7_75t_R n_4547 (.A1(n_4315_o_0),
    .A2(net59),
    .B(n_4258_o_0),
    .C(n_4314_o_0),
    .Y(n_4547_o_0));
 OAI31xp33_ASAP7_75t_R n_4548 (.A1(n_4258_o_0),
    .A2(n_4475_o_0),
    .A3(n_4546_o_0),
    .B(n_4547_o_0),
    .Y(n_4548_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4549 (.A1(n_2520_o_0),
    .A2(n_4272_o_0),
    .B(n_4544_o_0),
    .C(n_4548_o_0),
    .Y(n_4549_o_0));
 OA21x2_ASAP7_75t_R n_4550 (.A1(n_4542_o_0),
    .A2(n_4543_o_0),
    .B(n_4549_o_0),
    .Y(n_4550_o_0));
 OAI211xp5_ASAP7_75t_R n_4551 (.A1(net47),
    .A2(n_4290_o_0),
    .B(n_4354_o_0),
    .C(n_4317_o_0),
    .Y(n_4551_o_0));
 OAI21xp33_ASAP7_75t_R n_4552 (.A1(n_4258_o_0),
    .A2(n_4321_o_0),
    .B(n_4551_o_0),
    .Y(n_4552_o_0));
 NAND2xp33_ASAP7_75t_R n_4553 (.A(n_4226_o_0),
    .B(n_4244_o_0),
    .Y(n_4553_o_0));
 INVx1_ASAP7_75t_R n_4554 (.A(n_4553_o_0),
    .Y(n_4554_o_0));
 NOR3xp33_ASAP7_75t_R n_4555 (.A(n_4554_o_0),
    .B(n_4460_o_0),
    .C(n_4258_o_0),
    .Y(n_4555_o_0));
 AOI211xp5_ASAP7_75t_R n_4556 (.A1(n_4408_o_0),
    .A2(net47),
    .B(n_4329_o_0),
    .C(n_4447_o_0),
    .Y(n_4556_o_0));
 OAI31xp33_ASAP7_75t_R n_4557 (.A1(n_4307_o_0),
    .A2(n_4555_o_0),
    .A3(n_4556_o_0),
    .B(n_4305_o_0),
    .Y(n_4557_o_0));
 AOI21xp33_ASAP7_75t_R n_4558 (.A1(n_4307_o_0),
    .A2(n_4552_o_0),
    .B(n_4557_o_0),
    .Y(n_4558_o_0));
 AOI21xp33_ASAP7_75t_R n_4559 (.A1(n_4337_o_0),
    .A2(n_4550_o_0),
    .B(n_4558_o_0),
    .Y(n_4559_o_0));
 OAI21xp33_ASAP7_75t_R n_4560 (.A1(net59),
    .A2(net47),
    .B(n_4317_o_0),
    .Y(n_4560_o_0));
 OAI21xp33_ASAP7_75t_R n_4561 (.A1(net27),
    .A2(n_4242_o_0),
    .B(n_4560_o_0),
    .Y(n_4561_o_0));
 AOI31xp33_ASAP7_75t_R n_4562 (.A1(n_4258_o_0),
    .A2(n_4284_o_0),
    .A3(n_4314_o_0),
    .B(n_4278_o_0),
    .Y(n_4562_o_0));
 OAI31xp33_ASAP7_75t_R n_4563 (.A1(net62),
    .A2(net59),
    .A3(net27),
    .B(n_4562_o_0),
    .Y(n_4563_o_0));
 OAI21xp33_ASAP7_75t_R n_4564 (.A1(n_4274_o_0),
    .A2(n_4561_o_0),
    .B(n_4563_o_0),
    .Y(n_4564_o_0));
 NAND2xp33_ASAP7_75t_R n_4565 (.A(net47),
    .B(n_4431_o_0),
    .Y(n_4565_o_0));
 AOI21xp33_ASAP7_75t_R n_4566 (.A1(n_4565_o_0),
    .A2(n_4385_o_0),
    .B(n_4277_o_0),
    .Y(n_4566_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4567 (.A1(n_4383_o_0),
    .A2(net27),
    .B(n_4566_o_0),
    .C(n_4337_o_0),
    .Y(n_4567_o_0));
 OAI21xp33_ASAP7_75t_R n_4568 (.A1(n_4287_o_0),
    .A2(n_4244_o_0),
    .B(n_4317_o_0),
    .Y(n_4568_o_0));
 OA21x2_ASAP7_75t_R n_4569 (.A1(n_4355_o_0),
    .A2(n_4568_o_0),
    .B(n_4274_o_0),
    .Y(n_4569_o_0));
 OAI21xp33_ASAP7_75t_R n_4570 (.A1(n_4412_o_0),
    .A2(n_4506_o_0),
    .B(n_4569_o_0),
    .Y(n_4570_o_0));
 AOI21xp33_ASAP7_75t_R n_4571 (.A1(n_4567_o_0),
    .A2(n_4570_o_0),
    .B(n_4401_o_0),
    .Y(n_4571_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4572 (.A1(n_4305_o_0),
    .A2(n_4564_o_0),
    .B(n_4571_o_0),
    .C(n_4391_o_0),
    .Y(n_4572_o_0));
 OAI21xp33_ASAP7_75t_R n_4573 (.A1(n_4504_o_0),
    .A2(n_4559_o_0),
    .B(n_4572_o_0),
    .Y(n_4573_o_0));
 OAI21xp33_ASAP7_75t_R n_4574 (.A1(n_4528_o_0),
    .A2(n_4541_o_0),
    .B(n_4573_o_0),
    .Y(n_4574_o_0));
 OAI21xp33_ASAP7_75t_R n_4575 (.A1(n_4366_o_0),
    .A2(n_4508_o_0),
    .B(n_4278_o_0),
    .Y(n_4575_o_0));
 AOI21xp33_ASAP7_75t_R n_4576 (.A1(n_4385_o_0),
    .A2(n_4553_o_0),
    .B(n_4575_o_0),
    .Y(n_4576_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4577 (.A1(n_4406_o_0),
    .A2(n_4289_o_0),
    .B(n_4329_o_0),
    .C(n_4274_o_0),
    .Y(n_4577_o_0));
 AOI21xp33_ASAP7_75t_R n_4578 (.A1(n_4280_o_0),
    .A2(n_4553_o_0),
    .B(n_4577_o_0),
    .Y(n_4578_o_0));
 OAI21xp33_ASAP7_75t_R n_4579 (.A1(n_4576_o_0),
    .A2(n_4578_o_0),
    .B(n_4337_o_0),
    .Y(n_4579_o_0));
 INVx1_ASAP7_75t_R n_4580 (.A(n_4565_o_0),
    .Y(n_4580_o_0));
 NAND3xp33_ASAP7_75t_R n_4581 (.A(n_4377_o_0),
    .B(n_4553_o_0),
    .C(n_4263_o_0),
    .Y(n_4581_o_0));
 OAI31xp33_ASAP7_75t_R n_4582 (.A1(n_4330_o_0),
    .A2(n_4580_o_0),
    .A3(n_4329_o_0),
    .B(n_4581_o_0),
    .Y(n_4582_o_0));
 INVx1_ASAP7_75t_R n_4583 (.A(n_4380_o_0),
    .Y(n_4583_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4584 (.A1(n_4351_o_0),
    .A2(n_4315_o_0),
    .B(n_4258_o_0),
    .C(n_4274_o_0),
    .Y(n_4584_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4585 (.A1(n_4383_o_0),
    .A2(n_4583_o_0),
    .B(n_4584_o_0),
    .C(n_4464_o_0),
    .Y(n_4585_o_0));
 AO21x1_ASAP7_75t_R n_4586 (.A1(n_4278_o_0),
    .A2(n_4582_o_0),
    .B(n_4585_o_0),
    .Y(n_4586_o_0));
 NAND3xp33_ASAP7_75t_R n_4587 (.A(n_4579_o_0),
    .B(n_4586_o_0),
    .C(n_4346_o_0),
    .Y(n_4587_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4588 (.A1(n_4451_o_0),
    .A2(n_4367_o_0),
    .B(net27),
    .C(n_4284_o_0),
    .Y(n_4588_o_0));
 NAND3xp33_ASAP7_75t_R n_4589 (.A(n_4377_o_0),
    .B(n_4403_o_0),
    .C(n_4263_o_0),
    .Y(n_4589_o_0));
 OAI31xp33_ASAP7_75t_R n_4590 (.A1(n_4322_o_0),
    .A2(n_4546_o_0),
    .A3(n_4329_o_0),
    .B(n_4589_o_0),
    .Y(n_4590_o_0));
 AOI21xp33_ASAP7_75t_R n_4591 (.A1(n_4277_o_0),
    .A2(n_4590_o_0),
    .B(n_4464_o_0),
    .Y(n_4591_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4592 (.A1(n_4588_o_0),
    .A2(n_4274_o_0),
    .B(n_4591_o_0),
    .C(n_4346_o_0),
    .Y(n_4592_o_0));
 AOI21xp33_ASAP7_75t_R n_4593 (.A1(n_4241_o_0),
    .A2(n_4226_o_0),
    .B(n_4200_o_0),
    .Y(n_4593_o_0));
 OAI21xp33_ASAP7_75t_R n_4594 (.A1(n_4593_o_0),
    .A2(n_4361_o_0),
    .B(n_4274_o_0),
    .Y(n_4594_o_0));
 AOI21xp33_ASAP7_75t_R n_4595 (.A1(n_4368_o_0),
    .A2(n_4367_o_0),
    .B(n_4263_o_0),
    .Y(n_4595_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4596 (.A1(n_4283_o_0),
    .A2(n_4516_o_0),
    .B(n_4445_o_0),
    .C(n_4277_o_0),
    .Y(n_4596_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4597 (.A1(n_4495_o_0),
    .A2(n_4481_o_0),
    .B(n_4596_o_0),
    .C(n_4337_o_0),
    .Y(n_4597_o_0));
 OAI21xp33_ASAP7_75t_R n_4598 (.A1(n_4594_o_0),
    .A2(n_4595_o_0),
    .B(n_4597_o_0),
    .Y(n_4598_o_0));
 AOI21xp33_ASAP7_75t_R n_4599 (.A1(n_4592_o_0),
    .A2(n_4598_o_0),
    .B(n_4470_o_0),
    .Y(n_4599_o_0));
 OAI21xp33_ASAP7_75t_R n_4600 (.A1(n_4263_o_0),
    .A2(n_4351_o_0),
    .B(n_4521_o_0),
    .Y(n_4600_o_0));
 OA21x2_ASAP7_75t_R n_4601 (.A1(n_4546_o_0),
    .A2(n_4568_o_0),
    .B(n_4337_o_0),
    .Y(n_4601_o_0));
 OAI21xp33_ASAP7_75t_R n_4602 (.A1(n_4283_o_0),
    .A2(n_4361_o_0),
    .B(n_4601_o_0),
    .Y(n_4602_o_0));
 OAI21xp33_ASAP7_75t_R n_4603 (.A1(n_4304_o_0),
    .A2(n_4600_o_0),
    .B(n_4602_o_0),
    .Y(n_4603_o_0));
 NAND3xp33_ASAP7_75t_R n_4604 (.A(n_4289_o_0),
    .B(n_4263_o_0),
    .C(net62),
    .Y(n_4604_o_0));
 INVx1_ASAP7_75t_R n_4605 (.A(n_4604_o_0),
    .Y(n_4605_o_0));
 AOI21xp33_ASAP7_75t_R n_4606 (.A1(n_4289_o_0),
    .A2(n_4450_o_0),
    .B(n_4464_o_0),
    .Y(n_4606_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4607 (.A1(net62),
    .A2(net82),
    .B(n_4412_o_0),
    .C(n_4606_o_0),
    .Y(n_4607_o_0));
 OAI21xp33_ASAP7_75t_R n_4608 (.A1(n_4605_o_0),
    .A2(n_4304_o_0),
    .B(n_4607_o_0),
    .Y(n_4608_o_0));
 AOI22xp33_ASAP7_75t_R n_4609 (.A1(n_4603_o_0),
    .A2(n_4278_o_0),
    .B1(n_4413_o_0),
    .B2(n_4608_o_0),
    .Y(n_4609_o_0));
 OAI22xp33_ASAP7_75t_R n_4610 (.A1(n_4506_o_0),
    .A2(n_4412_o_0),
    .B1(n_4568_o_0),
    .B2(n_4593_o_0),
    .Y(n_4610_o_0));
 AOI21xp33_ASAP7_75t_R n_4611 (.A1(n_4278_o_0),
    .A2(n_4610_o_0),
    .B(n_4518_o_0),
    .Y(n_4611_o_0));
 NOR2xp33_ASAP7_75t_R n_4612 (.A(n_4290_o_0),
    .B(n_4292_o_0),
    .Y(n_4612_o_0));
 AO21x1_ASAP7_75t_R n_4613 (.A1(n_4351_o_0),
    .A2(n_4315_o_0),
    .B(n_4263_o_0),
    .Y(n_4613_o_0));
 OAI211xp5_ASAP7_75t_R n_4614 (.A1(n_4612_o_0),
    .A2(n_4361_o_0),
    .B(n_4613_o_0),
    .C(n_4277_o_0),
    .Y(n_4614_o_0));
 NAND2xp33_ASAP7_75t_R n_4615 (.A(n_4368_o_0),
    .B(n_4487_o_0),
    .Y(n_4615_o_0));
 INVx1_ASAP7_75t_R n_4616 (.A(n_4418_o_0),
    .Y(n_4616_o_0));
 AOI21xp33_ASAP7_75t_R n_4617 (.A1(n_4615_o_0),
    .A2(n_4616_o_0),
    .B(n_4304_o_0),
    .Y(n_4617_o_0));
 AOI21xp33_ASAP7_75t_R n_4618 (.A1(n_4614_o_0),
    .A2(n_4617_o_0),
    .B(n_4346_o_0),
    .Y(n_4618_o_0));
 OAI21xp33_ASAP7_75t_R n_4619 (.A1(n_4464_o_0),
    .A2(n_4611_o_0),
    .B(n_4618_o_0),
    .Y(n_4619_o_0));
 OAI21xp33_ASAP7_75t_R n_4620 (.A1(n_4391_o_0),
    .A2(n_4609_o_0),
    .B(n_4619_o_0),
    .Y(n_4620_o_0));
 AOI22xp33_ASAP7_75t_R n_4621 (.A1(n_4587_o_0),
    .A2(n_4599_o_0),
    .B1(n_4401_o_0),
    .B2(n_4620_o_0),
    .Y(n_4621_o_0));
 OAI22xp33_ASAP7_75t_R n_4622 (.A1(n_4355_o_0),
    .A2(n_4329_o_0),
    .B1(n_4258_o_0),
    .B2(n_4438_o_0),
    .Y(n_4622_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4623 (.A1(n_4475_o_0),
    .A2(n_4495_o_0),
    .B(n_4318_o_0),
    .C(n_4274_o_0),
    .Y(n_4623_o_0));
 AOI21xp33_ASAP7_75t_R n_4624 (.A1(n_4277_o_0),
    .A2(n_4622_o_0),
    .B(n_4623_o_0),
    .Y(n_4624_o_0));
 NOR2xp33_ASAP7_75t_R n_4625 (.A(n_4278_o_0),
    .B(n_4446_o_0),
    .Y(n_4625_o_0));
 AOI21xp33_ASAP7_75t_R n_4626 (.A1(n_4287_o_0),
    .A2(n_4263_o_0),
    .B(net47),
    .Y(n_4626_o_0));
 AOI211xp5_ASAP7_75t_R n_4627 (.A1(n_4546_o_0),
    .A2(n_4329_o_0),
    .B(n_4274_o_0),
    .C(n_4626_o_0),
    .Y(n_4627_o_0));
 OAI21xp33_ASAP7_75t_R n_4628 (.A1(n_4282_o_0),
    .A2(n_4241_o_0),
    .B(n_4200_o_0),
    .Y(n_4628_o_0));
 AOI211xp5_ASAP7_75t_R n_4629 (.A1(n_4327_o_0),
    .A2(n_4628_o_0),
    .B(n_4278_o_0),
    .C(n_4258_o_0),
    .Y(n_4629_o_0));
 NOR4xp25_ASAP7_75t_R n_4630 (.A(n_4625_o_0),
    .B(n_4627_o_0),
    .C(n_4629_o_0),
    .D(n_4464_o_0),
    .Y(n_4630_o_0));
 AOI21xp33_ASAP7_75t_R n_4631 (.A1(n_4305_o_0),
    .A2(n_4624_o_0),
    .B(n_4630_o_0),
    .Y(n_4631_o_0));
 OAI21xp33_ASAP7_75t_R n_4632 (.A1(n_4279_o_0),
    .A2(n_4473_o_0),
    .B(n_4278_o_0),
    .Y(n_4632_o_0));
 AOI211xp5_ASAP7_75t_R n_4633 (.A1(n_4280_o_0),
    .A2(n_4353_o_0),
    .B(n_4632_o_0),
    .C(n_4305_o_0),
    .Y(n_4633_o_0));
 INVx1_ASAP7_75t_R n_4634 (.A(n_4633_o_0),
    .Y(n_4634_o_0));
 NAND4xp25_ASAP7_75t_R n_4635 (.A(n_4326_o_0),
    .B(n_4404_o_0),
    .C(n_4305_o_0),
    .D(n_4274_o_0),
    .Y(n_4635_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4636 (.A1(n_4353_o_0),
    .A2(n_4280_o_0),
    .B(n_4632_o_0),
    .C(n_4635_o_0),
    .Y(n_4636_o_0));
 OAI21xp33_ASAP7_75t_R n_4637 (.A1(n_4508_o_0),
    .A2(n_4379_o_0),
    .B(n_4529_o_0),
    .Y(n_4637_o_0));
 INVx1_ASAP7_75t_R n_4638 (.A(n_4322_o_0),
    .Y(n_4638_o_0));
 OAI21xp33_ASAP7_75t_R n_4639 (.A1(n_4324_o_0),
    .A2(n_4313_o_0),
    .B(n_4638_o_0),
    .Y(n_4639_o_0));
 NOR3xp33_ASAP7_75t_R n_4640 (.A(n_4322_o_0),
    .B(n_4453_o_0),
    .C(n_4258_o_0),
    .Y(n_4640_o_0));
 INVx1_ASAP7_75t_R n_4641 (.A(n_4640_o_0),
    .Y(n_4641_o_0));
 OAI211xp5_ASAP7_75t_R n_4642 (.A1(n_4329_o_0),
    .A2(n_4639_o_0),
    .B(n_4641_o_0),
    .C(n_4274_o_0),
    .Y(n_4642_o_0));
 AOI21xp33_ASAP7_75t_R n_4643 (.A1(n_4637_o_0),
    .A2(n_4642_o_0),
    .B(n_4464_o_0),
    .Y(n_4643_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4644 (.A1(n_4634_o_0),
    .A2(n_4636_o_0),
    .B(n_4643_o_0),
    .C(n_4402_o_0),
    .Y(n_4644_o_0));
 OAI21xp33_ASAP7_75t_R n_4645 (.A1(n_4504_o_0),
    .A2(n_4631_o_0),
    .B(n_4644_o_0),
    .Y(n_4645_o_0));
 AOI21xp33_ASAP7_75t_R n_4646 (.A1(n_4463_o_0),
    .A2(n_4530_o_0),
    .B(n_4277_o_0),
    .Y(n_4646_o_0));
 OA21x2_ASAP7_75t_R n_4647 (.A1(n_4404_o_0),
    .A2(n_4407_o_0),
    .B(n_4646_o_0),
    .Y(n_4647_o_0));
 INVx1_ASAP7_75t_R n_4648 (.A(n_4432_o_0),
    .Y(n_4648_o_0));
 OAI211xp5_ASAP7_75t_R n_4649 (.A1(n_4289_o_0),
    .A2(n_4467_o_0),
    .B(n_4648_o_0),
    .C(n_4351_o_0),
    .Y(n_4649_o_0));
 OAI21xp33_ASAP7_75t_R n_4650 (.A1(n_4278_o_0),
    .A2(n_4649_o_0),
    .B(n_4305_o_0),
    .Y(n_4650_o_0));
 OAI21xp33_ASAP7_75t_R n_4651 (.A1(n_4647_o_0),
    .A2(n_4650_o_0),
    .B(n_4402_o_0),
    .Y(n_4651_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4652 (.A1(n_4382_o_0),
    .A2(n_4379_o_0),
    .B(n_4258_o_0),
    .C(n_4489_o_0),
    .Y(n_4652_o_0));
 NOR2xp33_ASAP7_75t_R n_4653 (.A(n_4258_o_0),
    .B(n_4475_o_0),
    .Y(n_4653_o_0));
 OAI21xp33_ASAP7_75t_R n_4654 (.A1(n_4407_o_0),
    .A2(n_4515_o_0),
    .B(n_4274_o_0),
    .Y(n_4654_o_0));
 AOI21xp33_ASAP7_75t_R n_4655 (.A1(n_4653_o_0),
    .A2(n_4545_o_0),
    .B(n_4654_o_0),
    .Y(n_4655_o_0));
 AOI311xp33_ASAP7_75t_R n_4656 (.A1(n_4490_o_0),
    .A2(n_4652_o_0),
    .A3(n_4278_o_0),
    .B(n_4305_o_0),
    .C(n_4655_o_0),
    .Y(n_4656_o_0));
 NAND3xp33_ASAP7_75t_R n_4657 (.A(n_4638_o_0),
    .B(n_4403_o_0),
    .C(net27),
    .Y(n_4657_o_0));
 OAI31xp33_ASAP7_75t_R n_4658 (.A1(net47),
    .A2(n_4258_o_0),
    .A3(n_4366_o_0),
    .B(n_4657_o_0),
    .Y(n_4658_o_0));
 OAI21xp33_ASAP7_75t_R n_4659 (.A1(n_4289_o_0),
    .A2(n_4467_o_0),
    .B(n_4307_o_0),
    .Y(n_4659_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4660 (.A1(n_4290_o_0),
    .A2(n_4329_o_0),
    .B(n_4659_o_0),
    .C(n_4305_o_0),
    .Y(n_4660_o_0));
 AOI21xp33_ASAP7_75t_R n_4661 (.A1(n_4277_o_0),
    .A2(n_4658_o_0),
    .B(n_4660_o_0),
    .Y(n_4661_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4662 (.A1(n_4593_o_0),
    .A2(n_4447_o_0),
    .B(net27),
    .C(n_4640_o_0),
    .Y(n_4662_o_0));
 INVx1_ASAP7_75t_R n_4663 (.A(n_4595_o_0),
    .Y(n_4663_o_0));
 AOI21xp33_ASAP7_75t_R n_4664 (.A1(n_4439_o_0),
    .A2(n_4663_o_0),
    .B(n_4277_o_0),
    .Y(n_4664_o_0));
 AOI211xp5_ASAP7_75t_R n_4665 (.A1(n_4274_o_0),
    .A2(n_4662_o_0),
    .B(n_4664_o_0),
    .C(n_4305_o_0),
    .Y(n_4665_o_0));
 OAI21xp33_ASAP7_75t_R n_4666 (.A1(n_4661_o_0),
    .A2(n_4665_o_0),
    .B(n_4401_o_0),
    .Y(n_4666_o_0));
 OAI211xp5_ASAP7_75t_R n_4667 (.A1(n_4651_o_0),
    .A2(n_4656_o_0),
    .B(n_4666_o_0),
    .C(n_4390_o_0),
    .Y(n_4667_o_0));
 OAI21xp33_ASAP7_75t_R n_4668 (.A1(n_4346_o_0),
    .A2(n_4645_o_0),
    .B(n_4667_o_0),
    .Y(n_4668_o_0));
 AOI22xp33_ASAP7_75t_R n_4669 (.A1(n_4501_o_0),
    .A2(n_4263_o_0),
    .B1(n_4411_o_0),
    .B2(net27),
    .Y(n_4669_o_0));
 NOR2xp33_ASAP7_75t_R n_4670 (.A(n_4337_o_0),
    .B(n_4568_o_0),
    .Y(n_4670_o_0));
 AOI31xp33_ASAP7_75t_R n_4671 (.A1(n_4263_o_0),
    .A2(n_4284_o_0),
    .A3(n_4501_o_0),
    .B(n_4670_o_0),
    .Y(n_4671_o_0));
 OAI21xp33_ASAP7_75t_R n_4672 (.A1(n_4305_o_0),
    .A2(n_4669_o_0),
    .B(n_4671_o_0),
    .Y(n_4672_o_0));
 OAI321xp33_ASAP7_75t_R n_4673 (.A1(n_4287_o_0),
    .A2(n_4282_o_0),
    .A3(n_4313_o_0),
    .B1(n_4360_o_0),
    .B2(net47),
    .C(n_4317_o_0),
    .Y(n_4673_o_0));
 OAI31xp33_ASAP7_75t_R n_4674 (.A1(n_4258_o_0),
    .A2(n_4460_o_0),
    .A3(n_4546_o_0),
    .B(n_4673_o_0),
    .Y(n_4674_o_0));
 AOI21xp33_ASAP7_75t_R n_4675 (.A1(n_4304_o_0),
    .A2(n_4674_o_0),
    .B(n_4307_o_0),
    .Y(n_4675_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4676 (.A1(n_4648_o_0),
    .A2(n_4293_o_0),
    .B(n_4337_o_0),
    .C(n_4675_o_0),
    .Y(n_4676_o_0));
 OAI21xp33_ASAP7_75t_R n_4677 (.A1(n_4277_o_0),
    .A2(n_4672_o_0),
    .B(n_4676_o_0),
    .Y(n_4677_o_0));
 NAND2xp33_ASAP7_75t_R n_4678 (.A(n_4244_o_0),
    .B(n_4317_o_0),
    .Y(n_4678_o_0));
 AOI31xp33_ASAP7_75t_R n_4679 (.A1(n_4263_o_0),
    .A2(n_4501_o_0),
    .A3(n_4545_o_0),
    .B(n_4464_o_0),
    .Y(n_4679_o_0));
 OAI31xp33_ASAP7_75t_R n_4680 (.A1(n_4258_o_0),
    .A2(n_4593_o_0),
    .A3(n_4322_o_0),
    .B(n_4305_o_0),
    .Y(n_4680_o_0));
 AOI21xp33_ASAP7_75t_R n_4681 (.A1(n_4385_o_0),
    .A2(n_4284_o_0),
    .B(n_4680_o_0),
    .Y(n_4681_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4682 (.A1(n_4678_o_0),
    .A2(n_4350_o_0),
    .B(n_4679_o_0),
    .C(n_4681_o_0),
    .Y(n_4682_o_0));
 NAND2xp33_ASAP7_75t_R n_4683 (.A(n_4317_o_0),
    .B(n_4241_o_0),
    .Y(n_4683_o_0));
 INVx1_ASAP7_75t_R n_4684 (.A(n_4368_o_0),
    .Y(n_4684_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4685 (.A1(n_4258_o_0),
    .A2(n_4447_o_0),
    .B(n_4683_o_0),
    .C(n_4684_o_0),
    .Y(n_4685_o_0));
 NAND3xp33_ASAP7_75t_R n_4686 (.A(n_4685_o_0),
    .B(n_4464_o_0),
    .C(n_4307_o_0),
    .Y(n_4686_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4687 (.A1(n_4318_o_0),
    .A2(n_4490_o_0),
    .B(n_4425_o_0),
    .C(n_4686_o_0),
    .Y(n_4687_o_0));
 AOI211xp5_ASAP7_75t_R n_4688 (.A1(n_4682_o_0),
    .A2(n_4277_o_0),
    .B(n_4390_o_0),
    .C(n_4687_o_0),
    .Y(n_4688_o_0));
 AOI21xp33_ASAP7_75t_R n_4689 (.A1(n_4346_o_0),
    .A2(n_4677_o_0),
    .B(n_4688_o_0),
    .Y(n_4689_o_0));
 NOR2xp33_ASAP7_75t_R n_4690 (.A(n_4612_o_0),
    .B(n_4259_o_0),
    .Y(n_4690_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4691 (.A1(n_4409_o_0),
    .A2(n_4553_o_0),
    .B(net27),
    .C(n_4307_o_0),
    .Y(n_4691_o_0));
 OAI211xp5_ASAP7_75t_R n_4692 (.A1(n_4292_o_0),
    .A2(net82),
    .B(n_4287_o_0),
    .C(n_4258_o_0),
    .Y(n_4692_o_0));
 INVx1_ASAP7_75t_R n_4693 (.A(n_4407_o_0),
    .Y(n_4693_o_0));
 AOI31xp33_ASAP7_75t_R n_4694 (.A1(n_4263_o_0),
    .A2(n_4693_o_0),
    .A3(n_4403_o_0),
    .B(n_4307_o_0),
    .Y(n_4694_o_0));
 AOI21xp33_ASAP7_75t_R n_4695 (.A1(n_4692_o_0),
    .A2(n_4694_o_0),
    .B(n_4304_o_0),
    .Y(n_4695_o_0));
 OAI21xp33_ASAP7_75t_R n_4696 (.A1(n_4690_o_0),
    .A2(n_4691_o_0),
    .B(n_4695_o_0),
    .Y(n_4696_o_0));
 NAND3xp33_ASAP7_75t_R n_4697 (.A(n_4613_o_0),
    .B(n_4307_o_0),
    .C(n_4361_o_0),
    .Y(n_4697_o_0));
 INVx1_ASAP7_75t_R n_4698 (.A(n_4653_o_0),
    .Y(n_4698_o_0));
 OAI211xp5_ASAP7_75t_R n_4699 (.A1(n_4366_o_0),
    .A2(n_4678_o_0),
    .B(n_4698_o_0),
    .C(n_4274_o_0),
    .Y(n_4699_o_0));
 NAND3xp33_ASAP7_75t_R n_4700 (.A(n_4697_o_0),
    .B(n_4699_o_0),
    .C(n_4337_o_0),
    .Y(n_4700_o_0));
 NOR2xp33_ASAP7_75t_R n_4701 (.A(n_4289_o_0),
    .B(n_4678_o_0),
    .Y(n_4701_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4702 (.A1(n_4462_o_0),
    .A2(n_4263_o_0),
    .B(n_4701_o_0),
    .C(n_4435_o_0),
    .Y(n_4702_o_0));
 OAI211xp5_ASAP7_75t_R n_4703 (.A1(n_4429_o_0),
    .A2(n_4438_o_0),
    .B(n_4517_o_0),
    .C(n_4278_o_0),
    .Y(n_4703_o_0));
 OAI21xp33_ASAP7_75t_R n_4704 (.A1(n_4278_o_0),
    .A2(n_4702_o_0),
    .B(n_4703_o_0),
    .Y(n_4704_o_0));
 NAND3xp33_ASAP7_75t_R n_4705 (.A(n_4454_o_0),
    .B(n_4315_o_0),
    .C(n_4263_o_0),
    .Y(n_4705_o_0));
 OAI31xp33_ASAP7_75t_R n_4706 (.A1(n_4593_o_0),
    .A2(n_4481_o_0),
    .A3(n_4329_o_0),
    .B(n_4705_o_0),
    .Y(n_4706_o_0));
 OAI21xp33_ASAP7_75t_R n_4707 (.A1(net59),
    .A2(n_4263_o_0),
    .B(n_4307_o_0),
    .Y(n_4707_o_0));
 OAI21xp33_ASAP7_75t_R n_4708 (.A1(n_4707_o_0),
    .A2(n_4640_o_0),
    .B(n_4305_o_0),
    .Y(n_4708_o_0));
 AOI21xp33_ASAP7_75t_R n_4709 (.A1(n_4277_o_0),
    .A2(n_4706_o_0),
    .B(n_4708_o_0),
    .Y(n_4709_o_0));
 AOI211xp5_ASAP7_75t_R n_4710 (.A1(n_4704_o_0),
    .A2(n_4304_o_0),
    .B(n_4345_o_0),
    .C(n_4709_o_0),
    .Y(n_4710_o_0));
 AOI311xp33_ASAP7_75t_R n_4711 (.A1(n_4345_o_0),
    .A2(n_4696_o_0),
    .A3(n_4700_o_0),
    .B(n_4401_o_0),
    .C(n_4710_o_0),
    .Y(n_4711_o_0));
 AO21x1_ASAP7_75t_R n_4712 (.A1(n_4689_o_0),
    .A2(n_4401_o_0),
    .B(n_4711_o_0),
    .Y(n_4712_o_0));
 AOI21xp33_ASAP7_75t_R n_4713 (.A1(net82),
    .A2(n_4367_o_0),
    .B(n_4263_o_0),
    .Y(n_4713_o_0));
 AOI21xp33_ASAP7_75t_R n_4714 (.A1(n_4329_o_0),
    .A2(n_4593_o_0),
    .B(n_4713_o_0),
    .Y(n_4714_o_0));
 AOI31xp33_ASAP7_75t_R n_4715 (.A1(n_4604_o_0),
    .A2(n_4561_o_0),
    .A3(n_4305_o_0),
    .B(n_4278_o_0),
    .Y(n_4715_o_0));
 OAI21xp33_ASAP7_75t_R n_4716 (.A1(n_4464_o_0),
    .A2(n_4714_o_0),
    .B(n_4715_o_0),
    .Y(n_4716_o_0));
 OAI21xp33_ASAP7_75t_R n_4717 (.A1(net47),
    .A2(n_4287_o_0),
    .B(n_4422_o_0),
    .Y(n_4717_o_0));
 OAI31xp33_ASAP7_75t_R n_4718 (.A1(n_4365_o_0),
    .A2(n_4407_o_0),
    .A3(n_4329_o_0),
    .B(n_4717_o_0),
    .Y(n_4718_o_0));
 INVx1_ASAP7_75t_R n_4719 (.A(n_4718_o_0),
    .Y(n_4719_o_0));
 NAND3xp33_ASAP7_75t_R n_4720 (.A(n_4462_o_0),
    .B(n_4377_o_0),
    .C(n_4263_o_0),
    .Y(n_4720_o_0));
 OAI31xp33_ASAP7_75t_R n_4721 (.A1(n_4321_o_0),
    .A2(n_4322_o_0),
    .A3(n_4329_o_0),
    .B(n_4720_o_0),
    .Y(n_4721_o_0));
 AOI21xp33_ASAP7_75t_R n_4722 (.A1(n_4464_o_0),
    .A2(n_4721_o_0),
    .B(n_4277_o_0),
    .Y(n_4722_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4723 (.A1(n_4305_o_0),
    .A2(n_4719_o_0),
    .B(n_4722_o_0),
    .C(n_4391_o_0),
    .Y(n_4723_o_0));
 OAI211xp5_ASAP7_75t_R n_4724 (.A1(n_4241_o_0),
    .A2(net62),
    .B(n_4351_o_0),
    .C(net27),
    .Y(n_4724_o_0));
 AOI21xp33_ASAP7_75t_R n_4725 (.A1(n_4530_o_0),
    .A2(n_4280_o_0),
    .B(n_4464_o_0),
    .Y(n_4725_o_0));
 AOI22xp33_ASAP7_75t_R n_4726 (.A1(n_4450_o_0),
    .A2(n_4408_o_0),
    .B1(n_4329_o_0),
    .B2(n_4382_o_0),
    .Y(n_4726_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4727 (.A1(n_4263_o_0),
    .A2(n_4351_o_0),
    .B(n_4726_o_0),
    .C(n_4304_o_0),
    .Y(n_4727_o_0));
 AOI211xp5_ASAP7_75t_R n_4728 (.A1(n_4724_o_0),
    .A2(n_4725_o_0),
    .B(n_4727_o_0),
    .C(n_4278_o_0),
    .Y(n_4728_o_0));
 AOI21xp33_ASAP7_75t_R n_4729 (.A1(n_4403_o_0),
    .A2(n_4463_o_0),
    .B(n_4464_o_0),
    .Y(n_4729_o_0));
 OAI21xp33_ASAP7_75t_R n_4730 (.A1(n_4678_o_0),
    .A2(n_4453_o_0),
    .B(n_4729_o_0),
    .Y(n_4730_o_0));
 AOI21xp33_ASAP7_75t_R n_4731 (.A1(net59),
    .A2(n_4263_o_0),
    .B(n_4304_o_0),
    .Y(n_4731_o_0));
 OAI21xp33_ASAP7_75t_R n_4732 (.A1(n_4366_o_0),
    .A2(n_4515_o_0),
    .B(n_4731_o_0),
    .Y(n_4732_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4733 (.A1(net27),
    .A2(n_4325_o_0),
    .B(n_4730_o_0),
    .C(n_4732_o_0),
    .D(n_4277_o_0),
    .Y(n_4733_o_0));
 NOR3xp33_ASAP7_75t_R n_4734 (.A(n_4728_o_0),
    .B(n_4733_o_0),
    .C(n_4390_o_0),
    .Y(n_4734_o_0));
 AOI21xp33_ASAP7_75t_R n_4735 (.A1(n_4716_o_0),
    .A2(n_4723_o_0),
    .B(n_4734_o_0),
    .Y(n_4735_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4736 (.A1(n_4368_o_0),
    .A2(net27),
    .B(n_4463_o_0),
    .C(n_4364_o_0),
    .Y(n_4736_o_0));
 OAI31xp33_ASAP7_75t_R n_4737 (.A1(n_4258_o_0),
    .A2(n_4321_o_0),
    .A3(n_4279_o_0),
    .B(n_4473_o_0),
    .Y(n_4737_o_0));
 AOI21xp33_ASAP7_75t_R n_4738 (.A1(n_4304_o_0),
    .A2(n_4737_o_0),
    .B(n_4307_o_0),
    .Y(n_4738_o_0));
 AOI21xp33_ASAP7_75t_R n_4739 (.A1(n_4315_o_0),
    .A2(n_4351_o_0),
    .B(n_4263_o_0),
    .Y(n_4739_o_0));
 AOI211xp5_ASAP7_75t_R n_4740 (.A1(n_4329_o_0),
    .A2(n_4460_o_0),
    .B(n_4739_o_0),
    .C(n_4305_o_0),
    .Y(n_4740_o_0));
 AOI211xp5_ASAP7_75t_R n_4741 (.A1(n_4683_o_0),
    .A2(net59),
    .B(n_4365_o_0),
    .C(n_4337_o_0),
    .Y(n_4741_o_0));
 OA21x2_ASAP7_75t_R n_4742 (.A1(n_4740_o_0),
    .A2(n_4741_o_0),
    .B(n_4307_o_0),
    .Y(n_4742_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4743 (.A1(n_4736_o_0),
    .A2(n_4337_o_0),
    .B(n_4738_o_0),
    .C(n_4742_o_0),
    .Y(n_4743_o_0));
 INVx1_ASAP7_75t_R n_4744 (.A(n_4543_o_0),
    .Y(n_4744_o_0));
 NOR3xp33_ASAP7_75t_R n_4745 (.A(n_4593_o_0),
    .B(n_4322_o_0),
    .C(n_4329_o_0),
    .Y(n_4745_o_0));
 INVx1_ASAP7_75t_R n_4746 (.A(n_4745_o_0),
    .Y(n_4746_o_0));
 AOI21xp33_ASAP7_75t_R n_4747 (.A1(n_4412_o_0),
    .A2(n_4746_o_0),
    .B(n_4278_o_0),
    .Y(n_4747_o_0));
 OAI21xp33_ASAP7_75t_R n_4748 (.A1(n_4744_o_0),
    .A2(n_4747_o_0),
    .B(n_4304_o_0),
    .Y(n_4748_o_0));
 OAI31xp33_ASAP7_75t_R n_4749 (.A1(n_4287_o_0),
    .A2(net27),
    .A3(net62),
    .B(n_4277_o_0),
    .Y(n_4749_o_0));
 NOR3xp33_ASAP7_75t_R n_4750 (.A(n_4546_o_0),
    .B(n_4460_o_0),
    .C(n_4329_o_0),
    .Y(n_4750_o_0));
 NAND2xp33_ASAP7_75t_R n_4751 (.A(net59),
    .B(net62),
    .Y(n_4751_o_0));
 NAND2xp33_ASAP7_75t_R n_4752 (.A(net82),
    .B(net47),
    .Y(n_4752_o_0));
 AOI31xp33_ASAP7_75t_R n_4753 (.A1(n_4263_o_0),
    .A2(n_4638_o_0),
    .A3(n_4403_o_0),
    .B(n_4277_o_0),
    .Y(n_4753_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4754 (.A1(n_4751_o_0),
    .A2(n_4752_o_0),
    .B(n_4329_o_0),
    .C(n_4753_o_0),
    .Y(n_4754_o_0));
 OAI211xp5_ASAP7_75t_R n_4755 (.A1(n_4749_o_0),
    .A2(n_4750_o_0),
    .B(n_4754_o_0),
    .C(n_4464_o_0),
    .Y(n_4755_o_0));
 AOI31xp33_ASAP7_75t_R n_4756 (.A1(n_4346_o_0),
    .A2(n_4748_o_0),
    .A3(n_4755_o_0),
    .B(n_4402_o_0),
    .Y(n_4756_o_0));
 OAI21xp33_ASAP7_75t_R n_4757 (.A1(n_4390_o_0),
    .A2(n_4743_o_0),
    .B(n_4756_o_0),
    .Y(n_4757_o_0));
 OAI21xp33_ASAP7_75t_R n_4758 (.A1(n_4470_o_0),
    .A2(n_4735_o_0),
    .B(n_4757_o_0),
    .Y(n_4758_o_0));
 INVx1_ASAP7_75t_R n_4759 (.A(n_4492_o_0),
    .Y(n_4759_o_0));
 OAI21xp33_ASAP7_75t_R n_4760 (.A1(n_4407_o_0),
    .A2(n_4264_o_0),
    .B(n_4305_o_0),
    .Y(n_4760_o_0));
 AOI21xp33_ASAP7_75t_R n_4761 (.A1(n_4327_o_0),
    .A2(n_4628_o_0),
    .B(n_4329_o_0),
    .Y(n_4761_o_0));
 AOI211xp5_ASAP7_75t_R n_4762 (.A1(n_4287_o_0),
    .A2(n_4450_o_0),
    .B(n_4760_o_0),
    .C(n_4761_o_0),
    .Y(n_4762_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4763 (.A1(n_4283_o_0),
    .A2(n_4361_o_0),
    .B(n_4759_o_0),
    .C(n_4762_o_0),
    .Y(n_4763_o_0));
 OAI31xp33_ASAP7_75t_R n_4764 (.A1(n_4304_o_0),
    .A2(n_4745_o_0),
    .A3(n_4463_o_0),
    .B(n_4307_o_0),
    .Y(n_4764_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4765 (.A1(net27),
    .A2(n_4536_o_0),
    .B(n_4729_o_0),
    .C(n_4537_o_0),
    .D(n_4764_o_0),
    .Y(n_4765_o_0));
 AOI21xp33_ASAP7_75t_R n_4766 (.A1(n_4277_o_0),
    .A2(n_4763_o_0),
    .B(n_4765_o_0),
    .Y(n_4766_o_0));
 AO21x1_ASAP7_75t_R n_4767 (.A1(n_4258_o_0),
    .A2(n_4481_o_0),
    .B(n_4425_o_0),
    .Y(n_4767_o_0));
 OA22x2_ASAP7_75t_R n_4768 (.A1(n_4473_o_0),
    .A2(n_4279_o_0),
    .B1(n_4258_o_0),
    .B2(n_4241_o_0),
    .Y(n_4768_o_0));
 AOI31xp33_ASAP7_75t_R n_4769 (.A1(n_4263_o_0),
    .A2(n_4354_o_0),
    .A3(n_4377_o_0),
    .B(n_4464_o_0),
    .Y(n_4769_o_0));
 OAI21xp33_ASAP7_75t_R n_4770 (.A1(n_4329_o_0),
    .A2(n_4407_o_0),
    .B(n_4769_o_0),
    .Y(n_4770_o_0));
 OAI21xp33_ASAP7_75t_R n_4771 (.A1(n_4304_o_0),
    .A2(n_4768_o_0),
    .B(n_4770_o_0),
    .Y(n_4771_o_0));
 AOI31xp33_ASAP7_75t_R n_4772 (.A1(n_4263_o_0),
    .A2(n_4638_o_0),
    .A3(n_4354_o_0),
    .B(n_4304_o_0),
    .Y(n_4772_o_0));
 AOI22xp33_ASAP7_75t_R n_4773 (.A1(n_4771_o_0),
    .A2(n_4274_o_0),
    .B1(n_4529_o_0),
    .B2(n_4772_o_0),
    .Y(n_4773_o_0));
 OAI211xp5_ASAP7_75t_R n_4774 (.A1(n_4767_o_0),
    .A2(n_4605_o_0),
    .B(n_4773_o_0),
    .C(n_4390_o_0),
    .Y(n_4774_o_0));
 OAI21xp33_ASAP7_75t_R n_4775 (.A1(n_4346_o_0),
    .A2(n_4766_o_0),
    .B(n_4774_o_0),
    .Y(n_4775_o_0));
 AO21x1_ASAP7_75t_R n_4776 (.A1(n_4530_o_0),
    .A2(n_4351_o_0),
    .B(net27),
    .Y(n_4776_o_0));
 OAI31xp33_ASAP7_75t_R n_4777 (.A1(net62),
    .A2(net82),
    .A3(n_4263_o_0),
    .B(n_4776_o_0),
    .Y(n_4777_o_0));
 OAI22xp33_ASAP7_75t_R n_4778 (.A1(n_4460_o_0),
    .A2(n_4380_o_0),
    .B1(n_4283_o_0),
    .B2(n_4322_o_0),
    .Y(n_4778_o_0));
 OAI21xp33_ASAP7_75t_R n_4779 (.A1(n_4257_o_0),
    .A2(n_4253_o_0),
    .B(n_4778_o_0),
    .Y(n_4779_o_0));
 NAND4xp25_ASAP7_75t_R n_4780 (.A(n_4530_o_0),
    .B(n_4377_o_0),
    .C(n_4317_o_0),
    .D(n_4258_o_0),
    .Y(n_4780_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4781 (.A1(n_4779_o_0),
    .A2(n_4780_o_0),
    .B(n_4278_o_0),
    .C(n_4337_o_0),
    .Y(n_4781_o_0));
 NOR3xp33_ASAP7_75t_R n_4782 (.A(n_4379_o_0),
    .B(n_4366_o_0),
    .C(n_4258_o_0),
    .Y(n_4782_o_0));
 OAI21xp33_ASAP7_75t_R n_4783 (.A1(n_4257_o_0),
    .A2(n_4253_o_0),
    .B(n_4244_o_0),
    .Y(n_4783_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4784 (.A1(n_4324_o_0),
    .A2(n_4783_o_0),
    .B(n_4329_o_0),
    .C(n_4290_o_0),
    .Y(n_4784_o_0));
 AOI22xp33_ASAP7_75t_R n_4785 (.A1(n_4782_o_0),
    .A2(n_4277_o_0),
    .B1(n_4307_o_0),
    .B2(n_4784_o_0),
    .Y(n_4785_o_0));
 OAI211xp5_ASAP7_75t_R n_4786 (.A1(n_4446_o_0),
    .A2(n_4278_o_0),
    .B(n_4785_o_0),
    .C(n_4305_o_0),
    .Y(n_4786_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4787 (.A1(n_4307_o_0),
    .A2(n_4777_o_0),
    .B(n_4781_o_0),
    .C(n_4786_o_0),
    .Y(n_4787_o_0));
 NAND2xp33_ASAP7_75t_R n_4788 (.A(n_4403_o_0),
    .B(n_4385_o_0),
    .Y(n_4788_o_0));
 OAI31xp33_ASAP7_75t_R n_4789 (.A1(n_4382_o_0),
    .A2(n_4554_o_0),
    .A3(n_4264_o_0),
    .B(n_4788_o_0),
    .Y(n_4789_o_0));
 OAI21xp33_ASAP7_75t_R n_4790 (.A1(n_4568_o_0),
    .A2(n_4593_o_0),
    .B(n_4274_o_0),
    .Y(n_4790_o_0));
 AOI21xp33_ASAP7_75t_R n_4791 (.A1(n_4454_o_0),
    .A2(n_4487_o_0),
    .B(n_4790_o_0),
    .Y(n_4791_o_0));
 AOI21xp33_ASAP7_75t_R n_4792 (.A1(n_4307_o_0),
    .A2(n_4789_o_0),
    .B(n_4791_o_0),
    .Y(n_4792_o_0));
 NOR2xp33_ASAP7_75t_R n_4793 (.A(n_4317_o_0),
    .B(n_4431_o_0),
    .Y(n_4793_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4794 (.A1(n_4451_o_0),
    .A2(n_4445_o_0),
    .B(n_4793_o_0),
    .C(n_4277_o_0),
    .Y(n_4794_o_0));
 NAND4xp25_ASAP7_75t_R n_4795 (.A(n_4263_o_0),
    .B(n_4287_o_0),
    .C(net47),
    .D(net59),
    .Y(n_4795_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4796 (.A1(n_4327_o_0),
    .A2(n_4628_o_0),
    .B(n_4329_o_0),
    .C(n_4795_o_0),
    .Y(n_4796_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4797 (.A1(n_4384_o_0),
    .A2(n_4796_o_0),
    .B(n_4307_o_0),
    .C(n_4464_o_0),
    .Y(n_4797_o_0));
 AOI21xp33_ASAP7_75t_R n_4798 (.A1(n_4794_o_0),
    .A2(n_4797_o_0),
    .B(n_4390_o_0),
    .Y(n_4798_o_0));
 OAI21xp33_ASAP7_75t_R n_4799 (.A1(n_4337_o_0),
    .A2(n_4792_o_0),
    .B(n_4798_o_0),
    .Y(n_4799_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4800 (.A1(n_4391_o_0),
    .A2(n_4787_o_0),
    .B(n_4799_o_0),
    .C(n_4470_o_0),
    .Y(n_4800_o_0));
 AO21x1_ASAP7_75t_R n_4801 (.A1(n_4775_o_0),
    .A2(n_4401_o_0),
    .B(n_4800_o_0),
    .Y(n_4801_o_0));
 XNOR2xp5_ASAP7_75t_R n_4802 (.A(_01024_),
    .B(_01032_),
    .Y(n_4802_o_0));
 INVx1_ASAP7_75t_R n_4803 (.A(n_4802_o_0),
    .Y(n_4803_o_0));
 XNOR2xp5_ASAP7_75t_R n_4804 (.A(_01073_),
    .B(_01112_),
    .Y(n_4804_o_0));
 XNOR2xp5_ASAP7_75t_R n_4805 (.A(_01033_),
    .B(n_4804_o_0),
    .Y(n_4805_o_0));
 NOR2xp33_ASAP7_75t_R n_4806 (.A(n_4803_o_0),
    .B(n_4805_o_0),
    .Y(n_4806_o_0));
 NOR2xp33_ASAP7_75t_R n_4807 (.A(_00711_),
    .B(net),
    .Y(n_4807_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4808 (.A1(n_4803_o_0),
    .A2(n_4805_o_0),
    .B(n_4806_o_0),
    .C(net),
    .D(n_4807_o_0),
    .Y(n_4808_o_0));
 NAND2xp33_ASAP7_75t_R n_4809 (.A(_00985_),
    .B(n_4808_o_0),
    .Y(n_4809_o_0));
 OAI21xp33_ASAP7_75t_R n_4810 (.A1(_00985_),
    .A2(n_4808_o_0),
    .B(n_4809_o_0),
    .Y(n_4810_o_0));
 INVx1_ASAP7_75t_R n_4811 (.A(n_4810_o_0),
    .Y(n_4811_o_0));
 XOR2xp5_ASAP7_75t_R n_4812 (.A(_01026_),
    .B(_01034_),
    .Y(n_4812_o_0));
 XNOR2xp5_ASAP7_75t_R n_4813 (.A(_01035_),
    .B(_01075_),
    .Y(n_4813_o_0));
 XNOR2xp5_ASAP7_75t_R n_4814 (.A(_01114_),
    .B(n_4813_o_0),
    .Y(n_4814_o_0));
 NAND2xp33_ASAP7_75t_R n_4815 (.A(n_4812_o_0),
    .B(n_4814_o_0),
    .Y(n_4815_o_0));
 OAI21xp33_ASAP7_75t_R n_4816 (.A1(n_4812_o_0),
    .A2(n_4814_o_0),
    .B(n_4815_o_0),
    .Y(n_4816_o_0));
 NOR2xp33_ASAP7_75t_R n_4817 (.A(_00709_),
    .B(net),
    .Y(n_4817_o_0));
 AOI211xp5_ASAP7_75t_R n_4818 (.A1(n_4816_o_0),
    .A2(net),
    .B(_00987_),
    .C(n_4817_o_0),
    .Y(n_4818_o_0));
 AOI21xp33_ASAP7_75t_R n_4819 (.A1(net),
    .A2(n_4816_o_0),
    .B(n_4817_o_0),
    .Y(n_4819_o_0));
 NOR2xp33_ASAP7_75t_R n_4820 (.A(n_2369_o_0),
    .B(n_4819_o_0),
    .Y(n_4820_o_0));
 NOR2xp33_ASAP7_75t_R n_4821 (.A(n_4818_o_0),
    .B(n_4820_o_0),
    .Y(n_4821_o_0));
 INVx1_ASAP7_75t_R n_4822 (.A(n_4821_o_0),
    .Y(n_4822_o_0));
 XOR2xp5_ASAP7_75t_R n_4823 (.A(_01025_),
    .B(_01033_),
    .Y(n_4823_o_0));
 XNOR2xp5_ASAP7_75t_R n_4824 (.A(_01034_),
    .B(_01074_),
    .Y(n_4824_o_0));
 XNOR2xp5_ASAP7_75t_R n_4825 (.A(_01113_),
    .B(n_4824_o_0),
    .Y(n_4825_o_0));
 NAND2xp33_ASAP7_75t_R n_4826 (.A(n_4823_o_0),
    .B(n_4825_o_0),
    .Y(n_4826_o_0));
 OAI21xp33_ASAP7_75t_R n_4827 (.A1(n_4823_o_0),
    .A2(n_4825_o_0),
    .B(n_4826_o_0),
    .Y(n_4827_o_0));
 NOR2xp33_ASAP7_75t_R n_4828 (.A(_00710_),
    .B(net),
    .Y(n_4828_o_0));
 AOI211xp5_ASAP7_75t_R n_4829 (.A1(n_4827_o_0),
    .A2(net),
    .B(n_2374_o_0),
    .C(n_4828_o_0),
    .Y(n_4829_o_0));
 AOI21xp33_ASAP7_75t_R n_4830 (.A1(net),
    .A2(n_4827_o_0),
    .B(n_4828_o_0),
    .Y(n_4830_o_0));
 NOR2xp33_ASAP7_75t_R n_4831 (.A(_00986_),
    .B(n_4830_o_0),
    .Y(n_4831_o_0));
 NOR2xp33_ASAP7_75t_R n_4832 (.A(n_4829_o_0),
    .B(n_4831_o_0),
    .Y(n_4832_o_0));
 INVx1_ASAP7_75t_R n_4833 (.A(_01031_),
    .Y(n_4833_o_0));
 XNOR2xp5_ASAP7_75t_R n_4834 (.A(_01022_),
    .B(_01027_),
    .Y(n_4834_o_0));
 XNOR2xp5_ASAP7_75t_R n_4835 (.A(n_4833_o_0),
    .B(n_4834_o_0),
    .Y(n_4835_o_0));
 XNOR2xp5_ASAP7_75t_R n_4836 (.A(_01030_),
    .B(_01035_),
    .Y(n_4836_o_0));
 XNOR2xp5_ASAP7_75t_R n_4837 (.A(_01071_),
    .B(_01110_),
    .Y(n_4837_o_0));
 XNOR2xp5_ASAP7_75t_R n_4838 (.A(n_4836_o_0),
    .B(n_4837_o_0),
    .Y(n_4838_o_0));
 XOR2xp5_ASAP7_75t_R n_4839 (.A(_01022_),
    .B(_01027_),
    .Y(n_4839_o_0));
 NAND2xp33_ASAP7_75t_R n_4840 (.A(n_4833_o_0),
    .B(n_4839_o_0),
    .Y(n_4840_o_0));
 NAND2xp33_ASAP7_75t_R n_4841 (.A(_01031_),
    .B(n_4834_o_0),
    .Y(n_4841_o_0));
 XOR2xp5_ASAP7_75t_R n_4842 (.A(_01071_),
    .B(_01110_),
    .Y(n_4842_o_0));
 NAND2xp33_ASAP7_75t_R n_4843 (.A(n_4836_o_0),
    .B(n_4842_o_0),
    .Y(n_4843_o_0));
 XOR2xp5_ASAP7_75t_R n_4844 (.A(_01030_),
    .B(_01035_),
    .Y(n_4844_o_0));
 NAND2xp33_ASAP7_75t_R n_4845 (.A(n_4837_o_0),
    .B(n_4844_o_0),
    .Y(n_4845_o_0));
 AOI22xp33_ASAP7_75t_R n_4846 (.A1(n_4840_o_0),
    .A2(n_4841_o_0),
    .B1(n_4843_o_0),
    .B2(n_4845_o_0),
    .Y(n_4846_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4847 (.A1(n_4835_o_0),
    .A2(n_4838_o_0),
    .B(n_4846_o_0),
    .C(net77),
    .Y(n_4847_o_0));
 OAI21xp33_ASAP7_75t_R n_4848 (.A1(_00713_),
    .A2(_00858_),
    .B(n_4847_o_0),
    .Y(n_4848_o_0));
 NOR2xp33_ASAP7_75t_R n_4849 (.A(n_4837_o_0),
    .B(n_4844_o_0),
    .Y(n_4849_o_0));
 NOR2xp33_ASAP7_75t_R n_4850 (.A(n_4836_o_0),
    .B(n_4842_o_0),
    .Y(n_4850_o_0));
 OAI21xp33_ASAP7_75t_R n_4851 (.A1(_01031_),
    .A2(n_4834_o_0),
    .B(n_4841_o_0),
    .Y(n_4851_o_0));
 NOR2xp33_ASAP7_75t_R n_4852 (.A(n_4833_o_0),
    .B(n_4839_o_0),
    .Y(n_4852_o_0));
 NOR2xp33_ASAP7_75t_R n_4853 (.A(_01031_),
    .B(n_4834_o_0),
    .Y(n_4853_o_0));
 OAI22xp33_ASAP7_75t_R n_4854 (.A1(n_4849_o_0),
    .A2(n_4850_o_0),
    .B1(n_4852_o_0),
    .B2(n_4853_o_0),
    .Y(n_4854_o_0));
 OAI31xp33_ASAP7_75t_R n_4855 (.A1(n_4849_o_0),
    .A2(n_4850_o_0),
    .A3(n_4851_o_0),
    .B(n_4854_o_0),
    .Y(n_4855_o_0));
 NOR2xp33_ASAP7_75t_R n_4856 (.A(_00713_),
    .B(net77),
    .Y(n_4856_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4857 (.A1(n_4855_o_0),
    .A2(net77),
    .B(n_4856_o_0),
    .C(_00983_),
    .Y(n_4857_o_0));
 OAI21x1_ASAP7_75t_R n_4858 (.A1(_00983_),
    .A2(n_4848_o_0),
    .B(n_4857_o_0),
    .Y(n_4858_o_0));
 INVx2_ASAP7_75t_R n_4859 (.A(n_4858_o_0),
    .Y(n_4859_o_0));
 NAND2xp33_ASAP7_75t_R n_4860 (.A(_01021_),
    .B(_01029_),
    .Y(n_4860_o_0));
 OAI21xp33_ASAP7_75t_R n_4861 (.A1(_01021_),
    .A2(_01029_),
    .B(n_4860_o_0),
    .Y(n_4861_o_0));
 INVx1_ASAP7_75t_R n_4862 (.A(n_4861_o_0),
    .Y(n_4862_o_0));
 XNOR2xp5_ASAP7_75t_R n_4863 (.A(_01070_),
    .B(_01109_),
    .Y(n_4863_o_0));
 XNOR2xp5_ASAP7_75t_R n_4864 (.A(_01030_),
    .B(n_4863_o_0),
    .Y(n_4864_o_0));
 INVx1_ASAP7_75t_R n_4865 (.A(_01070_),
    .Y(n_4865_o_0));
 NOR2xp33_ASAP7_75t_R n_4866 (.A(_01109_),
    .B(n_4865_o_0),
    .Y(n_4866_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4867 (.A1(n_4865_o_0),
    .A2(_01109_),
    .B(n_4866_o_0),
    .C(_01030_),
    .Y(n_4867_o_0));
 INVx1_ASAP7_75t_R n_4868 (.A(_01030_),
    .Y(n_4868_o_0));
 NAND2xp33_ASAP7_75t_R n_4869 (.A(n_4868_o_0),
    .B(n_4863_o_0),
    .Y(n_4869_o_0));
 AOI21xp33_ASAP7_75t_R n_4870 (.A1(n_4867_o_0),
    .A2(n_4869_o_0),
    .B(n_4862_o_0),
    .Y(n_4870_o_0));
 OAI21xp33_ASAP7_75t_R n_4871 (.A1(_00522_),
    .A2(net39),
    .B(n_2487_o_0),
    .Y(n_4871_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4872 (.A1(n_4862_o_0),
    .A2(n_4864_o_0),
    .B(n_4870_o_0),
    .C(net77),
    .D(n_4871_o_0),
    .Y(n_4872_o_0));
 INVx1_ASAP7_75t_R n_4873 (.A(n_4872_o_0),
    .Y(n_4873_o_0));
 INVx1_ASAP7_75t_R n_4874 (.A(_00522_),
    .Y(n_4874_o_0));
 NOR2xp33_ASAP7_75t_R n_4875 (.A(n_4868_o_0),
    .B(n_4863_o_0),
    .Y(n_4875_o_0));
 AOI211xp5_ASAP7_75t_R n_4876 (.A1(n_4863_o_0),
    .A2(n_4868_o_0),
    .B(n_4875_o_0),
    .C(n_4861_o_0),
    .Y(n_4876_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4877 (.A1(n_4869_o_0),
    .A2(n_4867_o_0),
    .B(n_4862_o_0),
    .C(net77),
    .Y(n_4877_o_0));
 OAI221xp5_ASAP7_75t_R n_4878 (.A1(n_4874_o_0),
    .A2(net),
    .B1(n_4876_o_0),
    .B2(n_4877_o_0),
    .C(_00982_),
    .Y(n_4878_o_0));
 XNOR2xp5_ASAP7_75t_R n_4879 (.A(_01027_),
    .B(_01035_),
    .Y(n_4879_o_0));
 INVx1_ASAP7_75t_R n_4880 (.A(_01107_),
    .Y(n_4880_o_0));
 INVx1_ASAP7_75t_R n_4881 (.A(_01035_),
    .Y(n_4881_o_0));
 NAND2xp33_ASAP7_75t_R n_4882 (.A(_01027_),
    .B(n_4881_o_0),
    .Y(n_4882_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4883 (.A1(n_4881_o_0),
    .A2(_01027_),
    .B(n_4882_o_0),
    .C(n_4880_o_0),
    .Y(n_4883_o_0));
 XNOR2xp5_ASAP7_75t_R n_4884 (.A(_01028_),
    .B(_01068_),
    .Y(n_4884_o_0));
 AOI211xp5_ASAP7_75t_R n_4885 (.A1(n_4879_o_0),
    .A2(n_4880_o_0),
    .B(n_4883_o_0),
    .C(n_4884_o_0),
    .Y(n_4885_o_0));
 NOR2xp33_ASAP7_75t_R n_4886 (.A(_01027_),
    .B(n_4881_o_0),
    .Y(n_4886_o_0));
 INVx1_ASAP7_75t_R n_4887 (.A(_01027_),
    .Y(n_4887_o_0));
 NOR2xp33_ASAP7_75t_R n_4888 (.A(_01035_),
    .B(n_4887_o_0),
    .Y(n_4888_o_0));
 OAI21xp33_ASAP7_75t_R n_4889 (.A1(n_4886_o_0),
    .A2(n_4888_o_0),
    .B(_01107_),
    .Y(n_4889_o_0));
 NAND2xp33_ASAP7_75t_R n_4890 (.A(n_4880_o_0),
    .B(n_4879_o_0),
    .Y(n_4890_o_0));
 XOR2xp5_ASAP7_75t_R n_4891 (.A(_01028_),
    .B(_01068_),
    .Y(n_4891_o_0));
 AOI21xp33_ASAP7_75t_R n_4892 (.A1(n_4889_o_0),
    .A2(n_4890_o_0),
    .B(n_4891_o_0),
    .Y(n_4892_o_0));
 NOR2xp33_ASAP7_75t_R n_4893 (.A(_00520_),
    .B(_00858_),
    .Y(n_4893_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4894 (.A1(n_4885_o_0),
    .A2(n_4892_o_0),
    .B(net39),
    .C(n_4893_o_0),
    .Y(n_4894_o_0));
 OAI311xp33_ASAP7_75t_R n_4895 (.A1(_01107_),
    .A2(n_4886_o_0),
    .A3(n_4888_o_0),
    .B1(n_4891_o_0),
    .C1(n_4889_o_0),
    .Y(n_4895_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4896 (.A1(n_4879_o_0),
    .A2(n_4880_o_0),
    .B(n_4883_o_0),
    .C(n_4884_o_0),
    .Y(n_4896_o_0));
 INVx1_ASAP7_75t_R n_4897 (.A(n_4893_o_0),
    .Y(n_4897_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4898 (.A1(n_4895_o_0),
    .A2(n_4896_o_0),
    .B(net5),
    .C(n_4897_o_0),
    .D(_00980_),
    .Y(n_4898_o_0));
 AOI21x1_ASAP7_75t_R n_4899 (.A1(_00980_),
    .A2(n_4894_o_0),
    .B(n_4898_o_0),
    .Y(n_4899_o_0));
 XNOR2xp5_ASAP7_75t_R n_4900 (.A(_01020_),
    .B(_01027_),
    .Y(n_4900_o_0));
 INVx1_ASAP7_75t_R n_4901 (.A(_01108_),
    .Y(n_4901_o_0));
 NAND2xp33_ASAP7_75t_R n_4902 (.A(_01020_),
    .B(n_4887_o_0),
    .Y(n_4902_o_0));
 OAI211xp5_ASAP7_75t_R n_4903 (.A1(n_4887_o_0),
    .A2(_01020_),
    .B(n_4902_o_0),
    .C(n_4901_o_0),
    .Y(n_4903_o_0));
 OAI21xp33_ASAP7_75t_R n_4904 (.A1(n_4900_o_0),
    .A2(n_4901_o_0),
    .B(n_4903_o_0),
    .Y(n_4904_o_0));
 NOR2xp33_ASAP7_75t_R n_4905 (.A(_01029_),
    .B(_01069_),
    .Y(n_4905_o_0));
 XNOR2xp5_ASAP7_75t_R n_4906 (.A(_01028_),
    .B(_01035_),
    .Y(n_4906_o_0));
 NAND2xp33_ASAP7_75t_R n_4907 (.A(_01029_),
    .B(_01069_),
    .Y(n_4907_o_0));
 INVx1_ASAP7_75t_R n_4908 (.A(n_4907_o_0),
    .Y(n_4908_o_0));
 NOR2xp33_ASAP7_75t_R n_4909 (.A(_01028_),
    .B(n_4881_o_0),
    .Y(n_4909_o_0));
 INVx1_ASAP7_75t_R n_4910 (.A(_01028_),
    .Y(n_4910_o_0));
 NOR2xp33_ASAP7_75t_R n_4911 (.A(_01035_),
    .B(n_4910_o_0),
    .Y(n_4911_o_0));
 XOR2xp5_ASAP7_75t_R n_4912 (.A(_01029_),
    .B(_01069_),
    .Y(n_4912_o_0));
 OAI33xp33_ASAP7_75t_R n_4913 (.A1(n_4905_o_0),
    .A2(n_4906_o_0),
    .A3(n_4908_o_0),
    .B1(n_4909_o_0),
    .B2(n_4911_o_0),
    .B3(n_4912_o_0),
    .Y(n_4913_o_0));
 NOR2xp33_ASAP7_75t_R n_4914 (.A(n_4901_o_0),
    .B(n_4900_o_0),
    .Y(n_4914_o_0));
 XOR2xp5_ASAP7_75t_R n_4915 (.A(_01020_),
    .B(_01027_),
    .Y(n_4915_o_0));
 NOR2xp33_ASAP7_75t_R n_4916 (.A(_01108_),
    .B(n_4915_o_0),
    .Y(n_4916_o_0));
 OAI21xp33_ASAP7_75t_R n_4917 (.A1(n_4914_o_0),
    .A2(n_4916_o_0),
    .B(n_4913_o_0),
    .Y(n_4917_o_0));
 OAI21xp33_ASAP7_75t_R n_4918 (.A1(n_4904_o_0),
    .A2(n_4913_o_0),
    .B(n_4917_o_0),
    .Y(n_4918_o_0));
 OAI21xp33_ASAP7_75t_R n_4919 (.A1(_00519_),
    .A2(net39),
    .B(_00981_),
    .Y(n_4919_o_0));
 INVx1_ASAP7_75t_R n_4920 (.A(_00519_),
    .Y(n_4920_o_0));
 NOR2xp33_ASAP7_75t_R n_4921 (.A(_01020_),
    .B(n_4887_o_0),
    .Y(n_4921_o_0));
 INVx1_ASAP7_75t_R n_4922 (.A(_01020_),
    .Y(n_4922_o_0));
 NOR2xp33_ASAP7_75t_R n_4923 (.A(_01027_),
    .B(n_4922_o_0),
    .Y(n_4923_o_0));
 OAI21xp33_ASAP7_75t_R n_4924 (.A1(n_4921_o_0),
    .A2(n_4923_o_0),
    .B(_01108_),
    .Y(n_4924_o_0));
 NAND2xp33_ASAP7_75t_R n_4925 (.A(_01028_),
    .B(n_4881_o_0),
    .Y(n_4925_o_0));
 OAI21xp33_ASAP7_75t_R n_4926 (.A1(_01029_),
    .A2(_01069_),
    .B(n_4907_o_0),
    .Y(n_4926_o_0));
 NAND2xp33_ASAP7_75t_R n_4927 (.A(_01035_),
    .B(n_4910_o_0),
    .Y(n_4927_o_0));
 XOR2xp5_ASAP7_75t_R n_4928 (.A(_01028_),
    .B(_01035_),
    .Y(n_4928_o_0));
 INVx1_ASAP7_75t_R n_4929 (.A(n_4905_o_0),
    .Y(n_4929_o_0));
 AOI33xp33_ASAP7_75t_R n_4930 (.A1(n_4925_o_0),
    .A2(n_4926_o_0),
    .A3(n_4927_o_0),
    .B1(n_4928_o_0),
    .B2(n_4929_o_0),
    .B3(n_4907_o_0),
    .Y(n_4930_o_0));
 AOI21xp33_ASAP7_75t_R n_4931 (.A1(n_4903_o_0),
    .A2(n_4924_o_0),
    .B(n_4930_o_0),
    .Y(n_4931_o_0));
 OAI31xp33_ASAP7_75t_R n_4932 (.A1(n_4916_o_0),
    .A2(n_4913_o_0),
    .A3(n_4914_o_0),
    .B(net77),
    .Y(n_4932_o_0));
 OAI221xp5_ASAP7_75t_R n_4933 (.A1(net39),
    .A2(n_4920_o_0),
    .B1(n_4931_o_0),
    .B2(n_4932_o_0),
    .C(n_2456_o_0),
    .Y(n_4933_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4934 (.A1(n_4918_o_0),
    .A2(net39),
    .B(n_4919_o_0),
    .C(n_4933_o_0),
    .Y(n_4934_o_0));
 NAND2xp33_ASAP7_75t_R n_4935 (.A(n_4899_o_0),
    .B(n_4934_o_0),
    .Y(n_4935_o_0));
 AOI21xp33_ASAP7_75t_R n_4936 (.A1(n_4873_o_0),
    .A2(n_4878_o_0),
    .B(n_4935_o_0),
    .Y(n_4936_o_0));
 OAI21xp33_ASAP7_75t_R n_4937 (.A1(n_4885_o_0),
    .A2(n_4892_o_0),
    .B(net),
    .Y(n_4937_o_0));
 OAI211xp5_ASAP7_75t_R n_4938 (.A1(_00520_),
    .A2(net),
    .B(n_4937_o_0),
    .C(_00980_),
    .Y(n_4938_o_0));
 XNOR2xp5_ASAP7_75t_R n_4939 (.A(_01108_),
    .B(n_4900_o_0),
    .Y(n_4939_o_0));
 OAI21xp33_ASAP7_75t_R n_4940 (.A1(n_4909_o_0),
    .A2(n_4911_o_0),
    .B(n_4912_o_0),
    .Y(n_4940_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4941 (.A1(_01029_),
    .A2(_01069_),
    .B(n_4905_o_0),
    .C(n_4906_o_0),
    .Y(n_4941_o_0));
 AOI22xp33_ASAP7_75t_R n_4942 (.A1(n_4940_o_0),
    .A2(n_4941_o_0),
    .B1(n_4924_o_0),
    .B2(n_4903_o_0),
    .Y(n_4942_o_0));
 AOI21xp33_ASAP7_75t_R n_4943 (.A1(n_4939_o_0),
    .A2(n_4930_o_0),
    .B(n_4942_o_0),
    .Y(n_4943_o_0));
 INVx1_ASAP7_75t_R n_4944 (.A(n_4919_o_0),
    .Y(n_4944_o_0));
 OAI21xp33_ASAP7_75t_R n_4945 (.A1(net2),
    .A2(n_4943_o_0),
    .B(n_4944_o_0),
    .Y(n_4945_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4946 (.A1(n_4890_o_0),
    .A2(n_4889_o_0),
    .B(n_4891_o_0),
    .C(n_4895_o_0),
    .Y(n_4946_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4947 (.A1(n_4946_o_0),
    .A2(net),
    .B(n_4893_o_0),
    .C(n_2432_o_0),
    .Y(n_4947_o_0));
 NAND4xp25_ASAP7_75t_R n_4948 (.A(n_4938_o_0),
    .B(n_4945_o_0),
    .C(n_4947_o_0),
    .D(n_4933_o_0),
    .Y(n_4948_o_0));
 AOI211xp5_ASAP7_75t_R n_4949 (.A1(n_4946_o_0),
    .A2(net),
    .B(n_2432_o_0),
    .C(n_4893_o_0),
    .Y(n_4949_o_0));
 OAI21xp33_ASAP7_75t_R n_4950 (.A1(n_4898_o_0),
    .A2(n_4949_o_0),
    .B(n_4934_o_0),
    .Y(n_4950_o_0));
 OA21x2_ASAP7_75t_R n_4951 (.A1(n_4877_o_0),
    .A2(n_4876_o_0),
    .B(_00982_),
    .Y(n_4951_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_4952 (.A1(n_4874_o_0),
    .A2(net39),
    .B(n_4951_o_0),
    .C(n_4872_o_0),
    .Y(n_4952_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4953 (.A1(n_4855_o_0),
    .A2(net39),
    .B(n_4856_o_0),
    .C(n_2411_o_0),
    .Y(n_4953_o_0));
 OAI21x1_ASAP7_75t_R n_4954 (.A1(n_4848_o_0),
    .A2(n_2411_o_0),
    .B(n_4953_o_0),
    .Y(n_4954_o_0));
 INVx1_ASAP7_75t_R n_4955 (.A(n_4954_o_0),
    .Y(n_4955_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4956 (.A1(n_4948_o_0),
    .A2(n_4950_o_0),
    .B(n_4952_o_0),
    .C(n_4955_o_0),
    .Y(n_4956_o_0));
 INVx1_ASAP7_75t_R n_4957 (.A(n_4956_o_0),
    .Y(n_4957_o_0));
 XNOR2xp5_ASAP7_75t_R n_4958 (.A(_01031_),
    .B(_01035_),
    .Y(n_4958_o_0));
 XNOR2xp5_ASAP7_75t_R n_4959 (.A(_01072_),
    .B(_01111_),
    .Y(n_4959_o_0));
 XNOR2xp5_ASAP7_75t_R n_4960 (.A(n_4958_o_0),
    .B(n_4959_o_0),
    .Y(n_4960_o_0));
 XNOR2xp5_ASAP7_75t_R n_4961 (.A(_01023_),
    .B(_01027_),
    .Y(n_4961_o_0));
 XOR2xp5_ASAP7_75t_R n_4962 (.A(_01032_),
    .B(n_4961_o_0),
    .Y(n_4962_o_0));
 AOI21xp33_ASAP7_75t_R n_4963 (.A1(n_4960_o_0),
    .A2(n_4962_o_0),
    .B(n_3021_o_0),
    .Y(n_4963_o_0));
 OA21x2_ASAP7_75t_R n_4964 (.A1(n_4960_o_0),
    .A2(n_4962_o_0),
    .B(n_4963_o_0),
    .Y(n_4964_o_0));
 AOI21xp33_ASAP7_75t_R n_4965 (.A1(net1),
    .A2(_00712_),
    .B(n_4964_o_0),
    .Y(n_4965_o_0));
 OR2x2_ASAP7_75t_R n_4966 (.A(_01032_),
    .B(n_4961_o_0),
    .Y(n_4966_o_0));
 NAND2xp33_ASAP7_75t_R n_4967 (.A(_01032_),
    .B(n_4961_o_0),
    .Y(n_4967_o_0));
 AO21x1_ASAP7_75t_R n_4968 (.A1(n_4966_o_0),
    .A2(n_4967_o_0),
    .B(n_4960_o_0),
    .Y(n_4968_o_0));
 AO221x1_ASAP7_75t_R n_4969 (.A1(_00712_),
    .A2(net9),
    .B1(n_4963_o_0),
    .B2(n_4968_o_0),
    .C(n_2521_o_0),
    .Y(n_4969_o_0));
 OAI21xp5_ASAP7_75t_R n_4970 (.A1(_00984_),
    .A2(n_4965_o_0),
    .B(n_4969_o_0),
    .Y(n_4970_o_0));
 NAND2xp33_ASAP7_75t_R n_4971 (.A(n_4913_o_0),
    .B(n_4904_o_0),
    .Y(n_4971_o_0));
 AOI21xp33_ASAP7_75t_R n_4972 (.A1(n_4930_o_0),
    .A2(n_4939_o_0),
    .B(net2),
    .Y(n_4972_o_0));
 AOI21xp33_ASAP7_75t_R n_4973 (.A1(n_4971_o_0),
    .A2(n_4972_o_0),
    .B(_00981_),
    .Y(n_4973_o_0));
 AOI21xp33_ASAP7_75t_R n_4974 (.A1(net77),
    .A2(n_4918_o_0),
    .B(n_4919_o_0),
    .Y(n_4974_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_4975 (.A1(n_4920_o_0),
    .A2(net),
    .B(n_4973_o_0),
    .C(n_4974_o_0),
    .Y(n_4975_o_0));
 AO21x1_ASAP7_75t_R n_4976 (.A1(n_4894_o_0),
    .A2(_00980_),
    .B(n_4898_o_0),
    .Y(n_4976_o_0));
 OA21x2_ASAP7_75t_R n_4977 (.A1(n_4877_o_0),
    .A2(n_4876_o_0),
    .B(_00982_),
    .Y(n_4977_o_0));
 OAI21xp33_ASAP7_75t_R n_4978 (.A1(_00522_),
    .A2(net),
    .B(n_2487_o_0),
    .Y(n_4978_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4979 (.A1(n_4862_o_0),
    .A2(n_4864_o_0),
    .B(n_4870_o_0),
    .C(net),
    .D(n_4978_o_0),
    .Y(n_4979_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4980 (.A1(n_4874_o_0),
    .A2(net),
    .B(n_4977_o_0),
    .C(n_4979_o_0),
    .Y(n_4980_o_0));
 NAND3xp33_ASAP7_75t_R n_4981 (.A(n_4975_o_0),
    .B(n_4976_o_0),
    .C(n_4980_o_0),
    .Y(n_4981_o_0));
 NOR2xp33_ASAP7_75t_R n_4982 (.A(n_4858_o_0),
    .B(n_4981_o_0),
    .Y(n_4982_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4983 (.A1(n_4859_o_0),
    .A2(n_4936_o_0),
    .B(n_4957_o_0),
    .C(n_4970_o_0),
    .D(n_4982_o_0),
    .Y(n_4983_o_0));
 AOI221xp5_ASAP7_75t_R n_4984 (.A1(net1),
    .A2(_00712_),
    .B1(n_4963_o_0),
    .B2(n_4968_o_0),
    .C(_00984_),
    .Y(n_4984_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_4985 (.A1(net9),
    .A2(_00712_),
    .B(n_4964_o_0),
    .C(_00984_),
    .D(n_4984_o_0),
    .Y(n_4985_o_0));
 INVx1_ASAP7_75t_R n_4986 (.A(n_4985_o_0),
    .Y(n_4986_o_0));
 OAI221xp5_ASAP7_75t_R n_4987 (.A1(n_4874_o_0),
    .A2(net),
    .B1(n_4876_o_0),
    .B2(n_4877_o_0),
    .C(_00982_),
    .Y(n_4987_o_0));
 INVx1_ASAP7_75t_R n_4988 (.A(n_4987_o_0),
    .Y(n_4988_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_4989 (.A1(n_4920_o_0),
    .A2(net),
    .B(n_4973_o_0),
    .C(n_4974_o_0),
    .Y(n_4989_o_0));
 OAI211xp5_ASAP7_75t_R n_4990 (.A1(n_4979_o_0),
    .A2(n_4988_o_0),
    .B(n_4989_o_0),
    .C(n_4899_o_0),
    .Y(n_4990_o_0));
 NAND2xp33_ASAP7_75t_R n_4991 (.A(n_4976_o_0),
    .B(n_4952_o_0),
    .Y(n_4991_o_0));
 NAND4xp25_ASAP7_75t_R n_4992 (.A(n_4986_o_0),
    .B(n_4990_o_0),
    .C(n_4991_o_0),
    .D(n_4858_o_0),
    .Y(n_4992_o_0));
 NAND2xp33_ASAP7_75t_R n_4993 (.A(n_4976_o_0),
    .B(n_4975_o_0),
    .Y(n_4993_o_0));
 OAI211xp5_ASAP7_75t_R n_4994 (.A1(n_4988_o_0),
    .A2(n_4979_o_0),
    .B(n_4945_o_0),
    .C(n_4933_o_0),
    .Y(n_4994_o_0));
 OAI21xp33_ASAP7_75t_R n_4995 (.A1(n_4899_o_0),
    .A2(n_4994_o_0),
    .B(n_4859_o_0),
    .Y(n_4995_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_4996 (.A1(n_4993_o_0),
    .A2(net60),
    .B(n_4995_o_0),
    .C(n_4986_o_0),
    .Y(n_4996_o_0));
 NAND2xp33_ASAP7_75t_R n_4997 (.A(n_4899_o_0),
    .B(n_4952_o_0),
    .Y(n_4997_o_0));
 NAND2xp5_ASAP7_75t_R n_4998 (.A(n_4878_o_0),
    .B(n_4873_o_0),
    .Y(n_4998_o_0));
 AOI221xp5_ASAP7_75t_R n_4999 (.A1(net9),
    .A2(_00519_),
    .B1(n_4971_o_0),
    .B2(n_4972_o_0),
    .C(_00981_),
    .Y(n_4999_o_0));
 OAI22xp33_ASAP7_75t_R n_5000 (.A1(n_4999_o_0),
    .A2(n_4974_o_0),
    .B1(n_4898_o_0),
    .B2(n_4949_o_0),
    .Y(n_5000_o_0));
 NAND2xp33_ASAP7_75t_R n_5001 (.A(n_4998_o_0),
    .B(n_5000_o_0),
    .Y(n_5001_o_0));
 INVx1_ASAP7_75t_R n_5002 (.A(n_4979_o_0),
    .Y(n_5002_o_0));
 NAND2xp33_ASAP7_75t_R n_5003 (.A(n_4987_o_0),
    .B(n_5002_o_0),
    .Y(n_5003_o_0));
 NOR2xp33_ASAP7_75t_R n_5004 (.A(n_5003_o_0),
    .B(n_5000_o_0),
    .Y(n_5004_o_0));
 NAND2xp33_ASAP7_75t_R n_5005 (.A(n_4859_o_0),
    .B(n_5004_o_0),
    .Y(n_5005_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5006 (.A1(n_4997_o_0),
    .A2(n_5001_o_0),
    .B(net95),
    .C(n_5005_o_0),
    .Y(n_5006_o_0));
 AOI21xp33_ASAP7_75t_R n_5007 (.A1(n_4933_o_0),
    .A2(n_4945_o_0),
    .B(n_4899_o_0),
    .Y(n_5007_o_0));
 AOI211xp5_ASAP7_75t_R n_5008 (.A1(n_4975_o_0),
    .A2(n_4899_o_0),
    .B(n_5007_o_0),
    .C(n_5003_o_0),
    .Y(n_5008_o_0));
 INVx1_ASAP7_75t_R n_5009 (.A(n_4970_o_0),
    .Y(n_5009_o_0));
 AOI21xp33_ASAP7_75t_R n_5010 (.A1(n_4859_o_0),
    .A2(n_5008_o_0),
    .B(n_5009_o_0),
    .Y(n_5010_o_0));
 OAI31xp33_ASAP7_75t_R n_5011 (.A1(net95),
    .A2(net60),
    .A3(net57),
    .B(n_5010_o_0),
    .Y(n_5011_o_0));
 OAI21xp33_ASAP7_75t_R n_5012 (.A1(n_4996_o_0),
    .A2(n_5006_o_0),
    .B(n_5011_o_0),
    .Y(n_5012_o_0));
 NAND2xp33_ASAP7_75t_R n_5013 (.A(n_2374_o_0),
    .B(n_4830_o_0),
    .Y(n_5013_o_0));
 OAI21xp33_ASAP7_75t_R n_5014 (.A1(n_4830_o_0),
    .A2(n_2374_o_0),
    .B(n_5013_o_0),
    .Y(n_5014_o_0));
 INVx1_ASAP7_75t_R n_5015 (.A(n_5014_o_0),
    .Y(n_5015_o_0));
 AOI32xp33_ASAP7_75t_R n_5016 (.A1(n_4832_o_0),
    .A2(n_4983_o_0),
    .A3(n_4992_o_0),
    .B1(n_5012_o_0),
    .B2(n_5015_o_0),
    .Y(n_5016_o_0));
 NAND2xp33_ASAP7_75t_R n_5017 (.A(n_4952_o_0),
    .B(n_4975_o_0),
    .Y(n_5017_o_0));
 INVx1_ASAP7_75t_R n_5018 (.A(n_5017_o_0),
    .Y(n_5018_o_0));
 INVx1_ASAP7_75t_R n_5019 (.A(n_4878_o_0),
    .Y(n_5019_o_0));
 OAI211xp5_ASAP7_75t_R n_5020 (.A1(n_4872_o_0),
    .A2(n_5019_o_0),
    .B(n_4948_o_0),
    .C(n_4950_o_0),
    .Y(n_5020_o_0));
 NAND2xp33_ASAP7_75t_R n_5021 (.A(net95),
    .B(n_5020_o_0),
    .Y(n_5021_o_0));
 OAI21xp33_ASAP7_75t_R n_5022 (.A1(n_4934_o_0),
    .A2(n_4976_o_0),
    .B(n_4950_o_0),
    .Y(n_5022_o_0));
 AOI21xp33_ASAP7_75t_R n_5023 (.A1(n_4952_o_0),
    .A2(n_5022_o_0),
    .B(n_4859_o_0),
    .Y(n_5023_o_0));
 INVx1_ASAP7_75t_R n_5024 (.A(n_5023_o_0),
    .Y(n_5024_o_0));
 OAI211xp5_ASAP7_75t_R n_5025 (.A1(n_5018_o_0),
    .A2(n_5021_o_0),
    .B(n_5024_o_0),
    .C(net51),
    .Y(n_5025_o_0));
 NAND2xp33_ASAP7_75t_R n_5026 (.A(n_4998_o_0),
    .B(n_4954_o_0),
    .Y(n_5026_o_0));
 INVx1_ASAP7_75t_R n_5027 (.A(n_5026_o_0),
    .Y(n_5027_o_0));
 NAND2xp33_ASAP7_75t_R n_5028 (.A(net60),
    .B(n_4954_o_0),
    .Y(n_5028_o_0));
 INVx1_ASAP7_75t_R n_5029 (.A(n_4935_o_0),
    .Y(n_5029_o_0));
 OAI22xp33_ASAP7_75t_R n_5030 (.A1(n_4956_o_0),
    .A2(n_5004_o_0),
    .B1(n_5028_o_0),
    .B2(n_5029_o_0),
    .Y(n_5030_o_0));
 AO21x1_ASAP7_75t_R n_5031 (.A1(n_5027_o_0),
    .A2(n_5000_o_0),
    .B(n_5030_o_0),
    .Y(n_5031_o_0));
 AOI21xp33_ASAP7_75t_R n_5032 (.A1(n_4986_o_0),
    .A2(n_5031_o_0),
    .B(n_5014_o_0),
    .Y(n_5032_o_0));
 NOR2xp33_ASAP7_75t_R n_5033 (.A(n_4952_o_0),
    .B(n_4975_o_0),
    .Y(n_5033_o_0));
 OAI21xp33_ASAP7_75t_R n_5034 (.A1(n_4934_o_0),
    .A2(n_4976_o_0),
    .B(n_4998_o_0),
    .Y(n_5034_o_0));
 NAND3xp33_ASAP7_75t_R n_5035 (.A(n_5034_o_0),
    .B(n_4991_o_0),
    .C(n_4858_o_0),
    .Y(n_5035_o_0));
 NOR2xp33_ASAP7_75t_R n_5036 (.A(net57),
    .B(n_4991_o_0),
    .Y(n_5036_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5037 (.A1(n_4955_o_0),
    .A2(n_5033_o_0),
    .B(n_5035_o_0),
    .C(n_5036_o_0),
    .Y(n_5037_o_0));
 NAND4xp25_ASAP7_75t_R n_5038 (.A(n_4986_o_0),
    .B(n_5001_o_0),
    .C(n_5017_o_0),
    .D(n_4954_o_0),
    .Y(n_5038_o_0));
 NAND3xp33_ASAP7_75t_R n_5039 (.A(n_4992_o_0),
    .B(n_5038_o_0),
    .C(n_4832_o_0),
    .Y(n_5039_o_0));
 NAND2xp33_ASAP7_75t_R n_5040 (.A(_00987_),
    .B(n_4819_o_0),
    .Y(n_5040_o_0));
 OAI21xp33_ASAP7_75t_R n_5041 (.A1(_00987_),
    .A2(n_4819_o_0),
    .B(n_5040_o_0),
    .Y(n_5041_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5042 (.A1(n_4970_o_0),
    .A2(n_5037_o_0),
    .B(n_5039_o_0),
    .C(n_5041_o_0),
    .Y(n_5042_o_0));
 AOI21xp33_ASAP7_75t_R n_5043 (.A1(n_5025_o_0),
    .A2(n_5032_o_0),
    .B(n_5042_o_0),
    .Y(n_5043_o_0));
 AOI21xp33_ASAP7_75t_R n_5044 (.A1(n_4822_o_0),
    .A2(n_5016_o_0),
    .B(n_5043_o_0),
    .Y(n_5044_o_0));
 NOR2xp33_ASAP7_75t_R n_5045 (.A(n_4952_o_0),
    .B(n_5000_o_0),
    .Y(n_5045_o_0));
 NOR2xp33_ASAP7_75t_R n_5046 (.A(n_4899_o_0),
    .B(n_4994_o_0),
    .Y(n_5046_o_0));
 NAND2xp33_ASAP7_75t_R n_5047 (.A(n_4952_o_0),
    .B(n_4935_o_0),
    .Y(n_5047_o_0));
 NAND2xp33_ASAP7_75t_R n_5048 (.A(n_4858_o_0),
    .B(n_5047_o_0),
    .Y(n_5048_o_0));
 OAI21xp33_ASAP7_75t_R n_5049 (.A1(n_5046_o_0),
    .A2(n_5048_o_0),
    .B(n_5009_o_0),
    .Y(n_5049_o_0));
 AOI21xp33_ASAP7_75t_R n_5050 (.A1(n_5045_o_0),
    .A2(net95),
    .B(n_5049_o_0),
    .Y(n_5050_o_0));
 NAND3xp33_ASAP7_75t_R n_5051 (.A(n_4980_o_0),
    .B(n_4934_o_0),
    .C(n_4899_o_0),
    .Y(n_5051_o_0));
 NAND2xp33_ASAP7_75t_R n_5052 (.A(n_4954_o_0),
    .B(n_5051_o_0),
    .Y(n_5052_o_0));
 AOI21xp33_ASAP7_75t_R n_5053 (.A1(n_4858_o_0),
    .A2(n_5045_o_0),
    .B(n_4986_o_0),
    .Y(n_5053_o_0));
 OA21x2_ASAP7_75t_R n_5054 (.A1(n_5052_o_0),
    .A2(n_5046_o_0),
    .B(n_5053_o_0),
    .Y(n_5054_o_0));
 AOI21xp33_ASAP7_75t_R n_5055 (.A1(n_4976_o_0),
    .A2(n_4975_o_0),
    .B(n_4952_o_0),
    .Y(n_5055_o_0));
 INVx1_ASAP7_75t_R n_5056 (.A(n_5055_o_0),
    .Y(n_5056_o_0));
 INVx1_ASAP7_75t_R n_5057 (.A(n_5001_o_0),
    .Y(n_5057_o_0));
 OAI31xp33_ASAP7_75t_R n_5058 (.A1(n_4955_o_0),
    .A2(n_5057_o_0),
    .A3(n_5004_o_0),
    .B(n_4985_o_0),
    .Y(n_5058_o_0));
 NOR2xp33_ASAP7_75t_R n_5059 (.A(n_4899_o_0),
    .B(n_4952_o_0),
    .Y(n_5059_o_0));
 INVx1_ASAP7_75t_R n_5060 (.A(n_5059_o_0),
    .Y(n_5060_o_0));
 NAND3xp33_ASAP7_75t_R n_5061 (.A(n_5060_o_0),
    .B(n_5051_o_0),
    .C(n_4858_o_0),
    .Y(n_5061_o_0));
 AOI211xp5_ASAP7_75t_R n_5062 (.A1(n_4873_o_0),
    .A2(n_4878_o_0),
    .B(n_4999_o_0),
    .C(n_4974_o_0),
    .Y(n_5062_o_0));
 INVx1_ASAP7_75t_R n_5063 (.A(n_5062_o_0),
    .Y(n_5063_o_0));
 NOR2xp33_ASAP7_75t_R n_5064 (.A(n_4955_o_0),
    .B(n_5008_o_0),
    .Y(n_5064_o_0));
 AOI21xp33_ASAP7_75t_R n_5065 (.A1(n_5063_o_0),
    .A2(n_5064_o_0),
    .B(n_4970_o_0),
    .Y(n_5065_o_0));
 AOI21xp33_ASAP7_75t_R n_5066 (.A1(n_5061_o_0),
    .A2(n_5065_o_0),
    .B(n_5015_o_0),
    .Y(n_5066_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5067 (.A1(n_4858_o_0),
    .A2(n_5056_o_0),
    .B(n_5058_o_0),
    .C(n_5066_o_0),
    .Y(n_5067_o_0));
 OAI31xp33_ASAP7_75t_R n_5068 (.A1(n_4832_o_0),
    .A2(n_5050_o_0),
    .A3(n_5054_o_0),
    .B(n_5067_o_0),
    .Y(n_5068_o_0));
 NOR3xp33_ASAP7_75t_R n_5069 (.A(n_5036_o_0),
    .B(n_5055_o_0),
    .C(n_4859_o_0),
    .Y(n_5069_o_0));
 NOR2xp67_ASAP7_75t_R n_5070 (.A(n_4899_o_0),
    .B(n_4998_o_0),
    .Y(n_5070_o_0));
 NOR2xp33_ASAP7_75t_R n_5071 (.A(n_4955_o_0),
    .B(n_5070_o_0),
    .Y(n_5071_o_0));
 OAI21xp33_ASAP7_75t_R n_5072 (.A1(net57),
    .A2(n_4991_o_0),
    .B(n_4954_o_0),
    .Y(n_5072_o_0));
 INVx1_ASAP7_75t_R n_5073 (.A(n_5072_o_0),
    .Y(n_5073_o_0));
 OAI21xp33_ASAP7_75t_R n_5074 (.A1(n_4934_o_0),
    .A2(n_4976_o_0),
    .B(n_4952_o_0),
    .Y(n_5074_o_0));
 NAND2xp33_ASAP7_75t_R n_5075 (.A(n_4858_o_0),
    .B(n_5074_o_0),
    .Y(n_5075_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5076 (.A1(n_4998_o_0),
    .A2(n_5022_o_0),
    .B(n_5075_o_0),
    .C(n_4985_o_0),
    .Y(n_5076_o_0));
 AO21x1_ASAP7_75t_R n_5077 (.A1(n_5073_o_0),
    .A2(n_5060_o_0),
    .B(n_5076_o_0),
    .Y(n_5077_o_0));
 OAI311xp33_ASAP7_75t_R n_5078 (.A1(n_4970_o_0),
    .A2(n_5069_o_0),
    .A3(n_5071_o_0),
    .B1(n_5014_o_0),
    .C1(n_5077_o_0),
    .Y(n_5078_o_0));
 OAI21xp33_ASAP7_75t_R n_5079 (.A1(n_4952_o_0),
    .A2(n_4976_o_0),
    .B(n_4954_o_0),
    .Y(n_5079_o_0));
 AOI21xp33_ASAP7_75t_R n_5080 (.A1(net57),
    .A2(n_4976_o_0),
    .B(n_5079_o_0),
    .Y(n_5080_o_0));
 NAND2xp33_ASAP7_75t_R n_5081 (.A(n_4976_o_0),
    .B(n_4975_o_0),
    .Y(n_5081_o_0));
 NAND3xp33_ASAP7_75t_R n_5082 (.A(n_5081_o_0),
    .B(n_4997_o_0),
    .C(n_4858_o_0),
    .Y(n_5082_o_0));
 INVx1_ASAP7_75t_R n_5083 (.A(n_5082_o_0),
    .Y(n_5083_o_0));
 INVx1_ASAP7_75t_R n_5084 (.A(n_4832_o_0),
    .Y(n_5084_o_0));
 NAND3xp33_ASAP7_75t_R n_5085 (.A(n_4975_o_0),
    .B(n_4899_o_0),
    .C(n_4952_o_0),
    .Y(n_5085_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5086 (.A1(n_4948_o_0),
    .A2(n_4950_o_0),
    .B(n_4952_o_0),
    .C(n_4859_o_0),
    .Y(n_5086_o_0));
 INVx1_ASAP7_75t_R n_5087 (.A(n_5086_o_0),
    .Y(n_5087_o_0));
 OAI31xp33_ASAP7_75t_R n_5088 (.A1(n_4859_o_0),
    .A2(n_5004_o_0),
    .A3(n_4936_o_0),
    .B(n_5009_o_0),
    .Y(n_5088_o_0));
 AO21x1_ASAP7_75t_R n_5089 (.A1(n_5085_o_0),
    .A2(n_5087_o_0),
    .B(n_5088_o_0),
    .Y(n_5089_o_0));
 OAI311xp33_ASAP7_75t_R n_5090 (.A1(n_4986_o_0),
    .A2(n_5080_o_0),
    .A3(n_5083_o_0),
    .B1(n_5084_o_0),
    .C1(n_5089_o_0),
    .Y(n_5090_o_0));
 NAND2xp33_ASAP7_75t_R n_5091 (.A(n_2393_o_0),
    .B(n_4808_o_0),
    .Y(n_5091_o_0));
 OAI21xp33_ASAP7_75t_R n_5092 (.A1(n_4808_o_0),
    .A2(n_2393_o_0),
    .B(n_5091_o_0),
    .Y(n_5092_o_0));
 INVx1_ASAP7_75t_R n_5093 (.A(n_5092_o_0),
    .Y(n_5093_o_0));
 AOI31xp33_ASAP7_75t_R n_5094 (.A1(n_5078_o_0),
    .A2(n_5090_o_0),
    .A3(n_4821_o_0),
    .B(n_5093_o_0),
    .Y(n_5094_o_0));
 OAI21xp33_ASAP7_75t_R n_5095 (.A1(n_5041_o_0),
    .A2(n_5068_o_0),
    .B(n_5094_o_0),
    .Y(n_5095_o_0));
 OAI21xp33_ASAP7_75t_R n_5096 (.A1(n_4811_o_0),
    .A2(n_5044_o_0),
    .B(n_5095_o_0),
    .Y(n_5096_o_0));
 AO21x1_ASAP7_75t_R n_5097 (.A1(n_5071_o_0),
    .A2(n_4990_o_0),
    .B(n_5092_o_0),
    .Y(n_5097_o_0));
 OAI211xp5_ASAP7_75t_R n_5098 (.A1(n_4952_o_0),
    .A2(n_4976_o_0),
    .B(n_4858_o_0),
    .C(net69),
    .Y(n_5098_o_0));
 OAI21xp33_ASAP7_75t_R n_5099 (.A1(n_5079_o_0),
    .A2(n_5004_o_0),
    .B(n_5098_o_0),
    .Y(n_5099_o_0));
 OAI22xp33_ASAP7_75t_R n_5100 (.A1(n_5097_o_0),
    .A2(n_4957_o_0),
    .B1(n_4810_o_0),
    .B2(n_5099_o_0),
    .Y(n_5100_o_0));
 NAND2xp33_ASAP7_75t_R n_5101 (.A(n_4934_o_0),
    .B(n_4952_o_0),
    .Y(n_5101_o_0));
 AND3x1_ASAP7_75t_R n_5102 (.A(n_4990_o_0),
    .B(n_5051_o_0),
    .C(n_4954_o_0),
    .Y(n_5102_o_0));
 AOI31xp33_ASAP7_75t_R n_5103 (.A1(n_4810_o_0),
    .A2(n_4858_o_0),
    .A3(n_5101_o_0),
    .B(n_5102_o_0),
    .Y(n_5103_o_0));
 AOI22xp33_ASAP7_75t_R n_5104 (.A1(n_5100_o_0),
    .A2(n_4832_o_0),
    .B1(n_5015_o_0),
    .B2(n_5103_o_0),
    .Y(n_5104_o_0));
 NOR2xp33_ASAP7_75t_R n_5105 (.A(n_4859_o_0),
    .B(n_5070_o_0),
    .Y(n_5105_o_0));
 NAND2xp33_ASAP7_75t_R n_5106 (.A(n_4899_o_0),
    .B(n_4934_o_0),
    .Y(n_5106_o_0));
 AO21x1_ASAP7_75t_R n_5107 (.A1(n_5105_o_0),
    .A2(n_5106_o_0),
    .B(n_5092_o_0),
    .Y(n_5107_o_0));
 AOI31xp33_ASAP7_75t_R n_5108 (.A1(n_4858_o_0),
    .A2(n_5020_o_0),
    .A3(n_5085_o_0),
    .B(n_4810_o_0),
    .Y(n_5108_o_0));
 OAI31xp33_ASAP7_75t_R n_5109 (.A1(n_4858_o_0),
    .A2(n_4993_o_0),
    .A3(net60),
    .B(n_5108_o_0),
    .Y(n_5109_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5110 (.A1(n_5060_o_0),
    .A2(n_5064_o_0),
    .B(n_5107_o_0),
    .C(n_5109_o_0),
    .Y(n_5110_o_0));
 AOI21xp33_ASAP7_75t_R n_5111 (.A1(net60),
    .A2(n_4993_o_0),
    .B(n_4995_o_0),
    .Y(n_5111_o_0));
 INVx1_ASAP7_75t_R n_5112 (.A(n_5034_o_0),
    .Y(n_5112_o_0));
 OAI21xp33_ASAP7_75t_R n_5113 (.A1(n_5112_o_0),
    .A2(n_5024_o_0),
    .B(n_5093_o_0),
    .Y(n_5113_o_0));
 AO21x1_ASAP7_75t_R n_5114 (.A1(n_5017_o_0),
    .A2(n_5106_o_0),
    .B(n_4858_o_0),
    .Y(n_5114_o_0));
 NAND2xp33_ASAP7_75t_R n_5115 (.A(n_4952_o_0),
    .B(n_4858_o_0),
    .Y(n_5115_o_0));
 INVx1_ASAP7_75t_R n_5116 (.A(n_5081_o_0),
    .Y(n_5116_o_0));
 OAI21xp33_ASAP7_75t_R n_5117 (.A1(n_5115_o_0),
    .A2(n_5116_o_0),
    .B(n_4811_o_0),
    .Y(n_5117_o_0));
 INVx1_ASAP7_75t_R n_5118 (.A(n_5117_o_0),
    .Y(n_5118_o_0));
 AOI21xp33_ASAP7_75t_R n_5119 (.A1(n_5114_o_0),
    .A2(n_5118_o_0),
    .B(n_4832_o_0),
    .Y(n_5119_o_0));
 OAI21xp33_ASAP7_75t_R n_5120 (.A1(n_5111_o_0),
    .A2(n_5113_o_0),
    .B(n_5119_o_0),
    .Y(n_5120_o_0));
 OAI21xp33_ASAP7_75t_R n_5121 (.A1(n_5110_o_0),
    .A2(n_5015_o_0),
    .B(n_5120_o_0),
    .Y(n_5121_o_0));
 OAI22xp33_ASAP7_75t_R n_5122 (.A1(n_4822_o_0),
    .A2(n_5104_o_0),
    .B1(n_5121_o_0),
    .B2(n_5041_o_0),
    .Y(n_5122_o_0));
 NOR2xp33_ASAP7_75t_R n_5123 (.A(n_4955_o_0),
    .B(n_5004_o_0),
    .Y(n_5123_o_0));
 AOI21xp33_ASAP7_75t_R n_5124 (.A1(n_5123_o_0),
    .A2(n_5060_o_0),
    .B(n_5117_o_0),
    .Y(n_5124_o_0));
 NAND2xp33_ASAP7_75t_R n_5125 (.A(n_4899_o_0),
    .B(n_4975_o_0),
    .Y(n_5125_o_0));
 NAND3xp33_ASAP7_75t_R n_5126 (.A(n_5125_o_0),
    .B(n_4858_o_0),
    .C(n_4998_o_0),
    .Y(n_5126_o_0));
 OA211x2_ASAP7_75t_R n_5127 (.A1(n_5018_o_0),
    .A2(n_5079_o_0),
    .B(n_5093_o_0),
    .C(n_5098_o_0),
    .Y(n_5127_o_0));
 AOI211xp5_ASAP7_75t_R n_5128 (.A1(n_5124_o_0),
    .A2(n_5126_o_0),
    .B(n_5127_o_0),
    .C(n_4832_o_0),
    .Y(n_5128_o_0));
 NAND2xp33_ASAP7_75t_R n_5129 (.A(n_4899_o_0),
    .B(net60),
    .Y(n_5129_o_0));
 NOR2xp33_ASAP7_75t_R n_5130 (.A(n_5129_o_0),
    .B(n_4955_o_0),
    .Y(n_5130_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5131 (.A1(n_5008_o_0),
    .A2(n_5057_o_0),
    .B(n_4955_o_0),
    .C(n_5130_o_0),
    .Y(n_5131_o_0));
 AOI21xp33_ASAP7_75t_R n_5132 (.A1(n_5045_o_0),
    .A2(net95),
    .B(n_4810_o_0),
    .Y(n_5132_o_0));
 AO21x1_ASAP7_75t_R n_5133 (.A1(n_5000_o_0),
    .A2(net60),
    .B(n_4858_o_0),
    .Y(n_5133_o_0));
 OAI21xp33_ASAP7_75t_R n_5134 (.A1(n_5112_o_0),
    .A2(n_5133_o_0),
    .B(n_5093_o_0),
    .Y(n_5134_o_0));
 AOI31xp33_ASAP7_75t_R n_5135 (.A1(n_4858_o_0),
    .A2(n_5020_o_0),
    .A3(n_5085_o_0),
    .B(n_5134_o_0),
    .Y(n_5135_o_0));
 AOI211xp5_ASAP7_75t_R n_5136 (.A1(n_5131_o_0),
    .A2(n_5132_o_0),
    .B(n_5135_o_0),
    .C(n_5015_o_0),
    .Y(n_5136_o_0));
 AOI31xp33_ASAP7_75t_R n_5137 (.A1(n_4976_o_0),
    .A2(n_4980_o_0),
    .A3(net69),
    .B(n_4956_o_0),
    .Y(n_5137_o_0));
 AOI31xp33_ASAP7_75t_R n_5138 (.A1(net95),
    .A2(n_4997_o_0),
    .A3(n_5001_o_0),
    .B(n_5137_o_0),
    .Y(n_5138_o_0));
 NOR2xp33_ASAP7_75t_R n_5139 (.A(n_4811_o_0),
    .B(n_5138_o_0),
    .Y(n_5139_o_0));
 NAND2xp33_ASAP7_75t_R n_5140 (.A(n_5125_o_0),
    .B(n_5027_o_0),
    .Y(n_5140_o_0));
 INVx1_ASAP7_75t_R n_5141 (.A(n_5074_o_0),
    .Y(n_5141_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5142 (.A1(n_4859_o_0),
    .A2(n_5033_o_0),
    .B(n_5140_o_0),
    .C(n_5141_o_0),
    .Y(n_5142_o_0));
 OAI21xp33_ASAP7_75t_R n_5143 (.A1(n_4810_o_0),
    .A2(n_5142_o_0),
    .B(n_5014_o_0),
    .Y(n_5143_o_0));
 AOI21xp33_ASAP7_75t_R n_5144 (.A1(net60),
    .A2(net69),
    .B(n_4954_o_0),
    .Y(n_5144_o_0));
 OR4x1_ASAP7_75t_R n_5145 (.A(n_4982_o_0),
    .B(n_5033_o_0),
    .C(n_5144_o_0),
    .D(n_4811_o_0),
    .Y(n_5145_o_0));
 AOI31xp33_ASAP7_75t_R n_5146 (.A1(n_4954_o_0),
    .A2(n_4997_o_0),
    .A3(n_5056_o_0),
    .B(n_4810_o_0),
    .Y(n_5146_o_0));
 OAI21xp33_ASAP7_75t_R n_5147 (.A1(n_5070_o_0),
    .A2(n_4956_o_0),
    .B(n_5146_o_0),
    .Y(n_5147_o_0));
 AOI31xp33_ASAP7_75t_R n_5148 (.A1(n_5015_o_0),
    .A2(n_5145_o_0),
    .A3(n_5147_o_0),
    .B(n_5041_o_0),
    .Y(n_5148_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5149 (.A1(n_5139_o_0),
    .A2(n_5143_o_0),
    .B(n_5148_o_0),
    .C(n_5009_o_0),
    .Y(n_5149_o_0));
 OAI31xp33_ASAP7_75t_R n_5150 (.A1(n_4822_o_0),
    .A2(n_5128_o_0),
    .A3(n_5136_o_0),
    .B(n_5149_o_0),
    .Y(n_5150_o_0));
 OAI21xp33_ASAP7_75t_R n_5151 (.A1(net51),
    .A2(n_5122_o_0),
    .B(n_5150_o_0),
    .Y(n_5151_o_0));
 OAI21xp33_ASAP7_75t_R n_5152 (.A1(n_5046_o_0),
    .A2(n_5024_o_0),
    .B(n_5009_o_0),
    .Y(n_5152_o_0));
 AOI31xp33_ASAP7_75t_R n_5153 (.A1(n_4998_o_0),
    .A2(net69),
    .A3(net95),
    .B(n_5152_o_0),
    .Y(n_5153_o_0));
 OAI21xp33_ASAP7_75t_R n_5154 (.A1(n_4975_o_0),
    .A2(n_4998_o_0),
    .B(n_4858_o_0),
    .Y(n_5154_o_0));
 OAI21xp33_ASAP7_75t_R n_5155 (.A1(n_5154_o_0),
    .A2(n_5059_o_0),
    .B(net51),
    .Y(n_5155_o_0));
 AOI21xp33_ASAP7_75t_R n_5156 (.A1(n_5064_o_0),
    .A2(n_5063_o_0),
    .B(n_5155_o_0),
    .Y(n_5156_o_0));
 AOI21xp33_ASAP7_75t_R n_5157 (.A1(n_4934_o_0),
    .A2(n_4976_o_0),
    .B(n_4998_o_0),
    .Y(n_5157_o_0));
 INVx1_ASAP7_75t_R n_5158 (.A(n_5157_o_0),
    .Y(n_5158_o_0));
 AOI22xp33_ASAP7_75t_R n_5159 (.A1(net57),
    .A2(n_4899_o_0),
    .B1(n_4873_o_0),
    .B2(n_4878_o_0),
    .Y(n_5159_o_0));
 NOR3xp33_ASAP7_75t_R n_5160 (.A(n_5008_o_0),
    .B(n_5159_o_0),
    .C(n_4859_o_0),
    .Y(n_5160_o_0));
 AOI31xp33_ASAP7_75t_R n_5161 (.A1(net95),
    .A2(n_5063_o_0),
    .A3(n_5158_o_0),
    .B(n_5160_o_0),
    .Y(n_5161_o_0));
 AOI21xp33_ASAP7_75t_R n_5162 (.A1(n_5106_o_0),
    .A2(n_5017_o_0),
    .B(n_4954_o_0),
    .Y(n_5162_o_0));
 AOI211xp5_ASAP7_75t_R n_5163 (.A1(net95),
    .A2(n_5101_o_0),
    .B(n_5162_o_0),
    .C(n_4970_o_0),
    .Y(n_5163_o_0));
 INVx1_ASAP7_75t_R n_5164 (.A(n_5163_o_0),
    .Y(n_5164_o_0));
 OAI211xp5_ASAP7_75t_R n_5165 (.A1(n_5161_o_0),
    .A2(n_5009_o_0),
    .B(n_5164_o_0),
    .C(n_5093_o_0),
    .Y(n_5165_o_0));
 OAI31xp33_ASAP7_75t_R n_5166 (.A1(n_5093_o_0),
    .A2(n_5153_o_0),
    .A3(n_5156_o_0),
    .B(n_5165_o_0),
    .Y(n_5166_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5167 (.A1(n_4873_o_0),
    .A2(n_4878_o_0),
    .B(n_4976_o_0),
    .C(n_4858_o_0),
    .Y(n_5167_o_0));
 INVx1_ASAP7_75t_R n_5168 (.A(n_5085_o_0),
    .Y(n_5168_o_0));
 OAI21xp33_ASAP7_75t_R n_5169 (.A1(n_5167_o_0),
    .A2(n_5168_o_0),
    .B(net51),
    .Y(n_5169_o_0));
 OAI21xp33_ASAP7_75t_R n_5170 (.A1(n_4934_o_0),
    .A2(n_4899_o_0),
    .B(n_4952_o_0),
    .Y(n_5170_o_0));
 AOI21xp33_ASAP7_75t_R n_5171 (.A1(n_5170_o_0),
    .A2(n_4957_o_0),
    .B(n_4970_o_0),
    .Y(n_5171_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5172 (.A1(net57),
    .A2(n_4976_o_0),
    .B(n_5026_o_0),
    .C(n_5171_o_0),
    .Y(n_5172_o_0));
 OAI211xp5_ASAP7_75t_R n_5173 (.A1(n_5169_o_0),
    .A2(n_5102_o_0),
    .B(n_5172_o_0),
    .C(n_5092_o_0),
    .Y(n_5173_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5174 (.A1(net69),
    .A2(n_4998_o_0),
    .B(n_4859_o_0),
    .C(n_5072_o_0),
    .Y(n_5174_o_0));
 NAND2xp33_ASAP7_75t_R n_5175 (.A(n_4975_o_0),
    .B(n_5070_o_0),
    .Y(n_5175_o_0));
 AOI31xp33_ASAP7_75t_R n_5176 (.A1(n_4955_o_0),
    .A2(n_5175_o_0),
    .A3(n_4994_o_0),
    .B(n_4986_o_0),
    .Y(n_5176_o_0));
 OAI31xp33_ASAP7_75t_R n_5177 (.A1(n_4998_o_0),
    .A2(net57),
    .A3(n_4955_o_0),
    .B(n_5176_o_0),
    .Y(n_5177_o_0));
 OAI211xp5_ASAP7_75t_R n_5178 (.A1(n_4970_o_0),
    .A2(n_5174_o_0),
    .B(n_5177_o_0),
    .C(n_4810_o_0),
    .Y(n_5178_o_0));
 AOI21xp33_ASAP7_75t_R n_5179 (.A1(n_5173_o_0),
    .A2(n_5178_o_0),
    .B(n_4832_o_0),
    .Y(n_5179_o_0));
 AOI21xp33_ASAP7_75t_R n_5180 (.A1(n_5014_o_0),
    .A2(n_5166_o_0),
    .B(n_5179_o_0),
    .Y(n_5180_o_0));
 NOR2xp33_ASAP7_75t_R n_5181 (.A(n_4976_o_0),
    .B(n_4952_o_0),
    .Y(n_5181_o_0));
 NAND2xp33_ASAP7_75t_R n_5182 (.A(n_4934_o_0),
    .B(n_4952_o_0),
    .Y(n_5182_o_0));
 NAND3xp33_ASAP7_75t_R n_5183 (.A(n_5020_o_0),
    .B(n_5182_o_0),
    .C(n_4954_o_0),
    .Y(n_5183_o_0));
 OAI31xp33_ASAP7_75t_R n_5184 (.A1(n_4859_o_0),
    .A2(n_5004_o_0),
    .A3(n_5181_o_0),
    .B(n_5183_o_0),
    .Y(n_5184_o_0));
 NOR3xp33_ASAP7_75t_R n_5185 (.A(n_5168_o_0),
    .B(n_5112_o_0),
    .C(n_4859_o_0),
    .Y(n_5185_o_0));
 NOR4xp25_ASAP7_75t_R n_5186 (.A(n_5185_o_0),
    .B(n_4970_o_0),
    .C(n_4810_o_0),
    .D(n_5073_o_0),
    .Y(n_5186_o_0));
 OAI211xp5_ASAP7_75t_R n_5187 (.A1(n_4991_o_0),
    .A2(net57),
    .B(n_4955_o_0),
    .C(n_4994_o_0),
    .Y(n_5187_o_0));
 OAI31xp33_ASAP7_75t_R n_5188 (.A1(n_4955_o_0),
    .A2(n_5055_o_0),
    .A3(n_5141_o_0),
    .B(n_5187_o_0),
    .Y(n_5188_o_0));
 NAND3xp33_ASAP7_75t_R n_5189 (.A(n_4948_o_0),
    .B(n_4950_o_0),
    .C(n_4980_o_0),
    .Y(n_5189_o_0));
 NAND2xp33_ASAP7_75t_R n_5190 (.A(n_4954_o_0),
    .B(n_5189_o_0),
    .Y(n_5190_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5191 (.A1(n_5062_o_0),
    .A2(n_5190_o_0),
    .B(n_5009_o_0),
    .C(n_4810_o_0),
    .Y(n_5191_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5192 (.A1(n_4899_o_0),
    .A2(n_4994_o_0),
    .B(n_5170_o_0),
    .C(n_4954_o_0),
    .Y(n_5192_o_0));
 AOI221xp5_ASAP7_75t_R n_5193 (.A1(n_4810_o_0),
    .A2(n_5192_o_0),
    .B1(n_5063_o_0),
    .B2(n_5064_o_0),
    .C(n_4970_o_0),
    .Y(n_5193_o_0));
 AOI211xp5_ASAP7_75t_R n_5194 (.A1(n_4970_o_0),
    .A2(n_5188_o_0),
    .B(n_5191_o_0),
    .C(n_5193_o_0),
    .Y(n_5194_o_0));
 AOI311xp33_ASAP7_75t_R n_5195 (.A1(n_4970_o_0),
    .A2(n_5092_o_0),
    .A3(n_5184_o_0),
    .B(n_5186_o_0),
    .C(n_5194_o_0),
    .Y(n_5195_o_0));
 INVx1_ASAP7_75t_R n_5196 (.A(n_5181_o_0),
    .Y(n_5196_o_0));
 OAI31xp33_ASAP7_75t_R n_5197 (.A1(n_4976_o_0),
    .A2(n_4998_o_0),
    .A3(n_4934_o_0),
    .B(n_4954_o_0),
    .Y(n_5197_o_0));
 AOI22xp33_ASAP7_75t_R n_5198 (.A1(n_4936_o_0),
    .A2(n_4859_o_0),
    .B1(n_4985_o_0),
    .B2(n_5197_o_0),
    .Y(n_5198_o_0));
 AOI31xp33_ASAP7_75t_R n_5199 (.A1(n_4858_o_0),
    .A2(n_4981_o_0),
    .A3(n_5196_o_0),
    .B(n_5198_o_0),
    .Y(n_5199_o_0));
 INVx1_ASAP7_75t_R n_5200 (.A(n_5170_o_0),
    .Y(n_5200_o_0));
 AOI21xp33_ASAP7_75t_R n_5201 (.A1(net69),
    .A2(n_4858_o_0),
    .B(net60),
    .Y(n_5201_o_0));
 NOR3xp33_ASAP7_75t_R n_5202 (.A(n_5200_o_0),
    .B(n_5201_o_0),
    .C(net51),
    .Y(n_5202_o_0));
 INVx1_ASAP7_75t_R n_5203 (.A(n_5182_o_0),
    .Y(n_5203_o_0));
 NOR4xp25_ASAP7_75t_R n_5204 (.A(n_5093_o_0),
    .B(n_5203_o_0),
    .C(n_4859_o_0),
    .D(n_4936_o_0),
    .Y(n_5204_o_0));
 OA21x2_ASAP7_75t_R n_5205 (.A1(n_5181_o_0),
    .A2(n_5197_o_0),
    .B(n_4985_o_0),
    .Y(n_5205_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5206 (.A1(n_5197_o_0),
    .A2(n_5181_o_0),
    .B(n_4985_o_0),
    .C(n_5093_o_0),
    .Y(n_5206_o_0));
 INVx1_ASAP7_75t_R n_5207 (.A(n_5020_o_0),
    .Y(n_5207_o_0));
 INVx1_ASAP7_75t_R n_5208 (.A(n_5079_o_0),
    .Y(n_5208_o_0));
 AOI21xp33_ASAP7_75t_R n_5209 (.A1(n_5051_o_0),
    .A2(n_5208_o_0),
    .B(n_4970_o_0),
    .Y(n_5209_o_0));
 OAI21xp33_ASAP7_75t_R n_5210 (.A1(n_5207_o_0),
    .A2(n_5024_o_0),
    .B(n_5209_o_0),
    .Y(n_5210_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5211 (.A1(n_5204_o_0),
    .A2(n_5205_o_0),
    .B(n_5206_o_0),
    .C(n_5210_o_0),
    .Y(n_5211_o_0));
 OAI311xp33_ASAP7_75t_R n_5212 (.A1(n_4811_o_0),
    .A2(n_5199_o_0),
    .A3(n_5202_o_0),
    .B1(n_4832_o_0),
    .C1(n_5211_o_0),
    .Y(n_5212_o_0));
 INVx1_ASAP7_75t_R n_5213 (.A(n_5212_o_0),
    .Y(n_5213_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5214 (.A1(n_5195_o_0),
    .A2(n_5084_o_0),
    .B(n_5213_o_0),
    .C(n_5041_o_0),
    .Y(n_5214_o_0));
 OAI21xp33_ASAP7_75t_R n_5215 (.A1(n_4821_o_0),
    .A2(n_5180_o_0),
    .B(n_5214_o_0),
    .Y(n_5215_o_0));
 INVx1_ASAP7_75t_R n_5216 (.A(n_4997_o_0),
    .Y(n_5216_o_0));
 OAI31xp33_ASAP7_75t_R n_5217 (.A1(n_4955_o_0),
    .A2(n_5216_o_0),
    .A3(n_5159_o_0),
    .B(net51),
    .Y(n_5217_o_0));
 OAI31xp33_ASAP7_75t_R n_5218 (.A1(n_4859_o_0),
    .A2(n_5112_o_0),
    .A3(n_5200_o_0),
    .B(n_5183_o_0),
    .Y(n_5218_o_0));
 AOI21xp33_ASAP7_75t_R n_5219 (.A1(n_4986_o_0),
    .A2(n_5218_o_0),
    .B(n_4810_o_0),
    .Y(n_5219_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5220 (.A1(n_5001_o_0),
    .A2(n_5023_o_0),
    .B(n_5217_o_0),
    .C(n_5219_o_0),
    .Y(n_5220_o_0));
 AOI31xp33_ASAP7_75t_R n_5221 (.A1(net95),
    .A2(n_5060_o_0),
    .A3(n_5182_o_0),
    .B(n_5023_o_0),
    .Y(n_5221_o_0));
 OAI21xp33_ASAP7_75t_R n_5222 (.A1(n_4956_o_0),
    .A2(n_5203_o_0),
    .B(n_5009_o_0),
    .Y(n_5222_o_0));
 AOI21xp33_ASAP7_75t_R n_5223 (.A1(n_5208_o_0),
    .A2(n_5081_o_0),
    .B(n_5222_o_0),
    .Y(n_5223_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5224 (.A1(net51),
    .A2(n_5221_o_0),
    .B(n_5223_o_0),
    .C(n_5093_o_0),
    .Y(n_5224_o_0));
 AOI21xp33_ASAP7_75t_R n_5225 (.A1(n_5081_o_0),
    .A2(n_5196_o_0),
    .B(n_4858_o_0),
    .Y(n_5225_o_0));
 NAND2xp33_ASAP7_75t_R n_5226 (.A(n_4986_o_0),
    .B(n_5175_o_0),
    .Y(n_5226_o_0));
 NAND3xp33_ASAP7_75t_R n_5227 (.A(n_5047_o_0),
    .B(n_5020_o_0),
    .C(net95),
    .Y(n_5227_o_0));
 OAI31xp33_ASAP7_75t_R n_5228 (.A1(n_4859_o_0),
    .A2(n_5033_o_0),
    .A3(n_5141_o_0),
    .B(n_5227_o_0),
    .Y(n_5228_o_0));
 AOI21xp33_ASAP7_75t_R n_5229 (.A1(n_4970_o_0),
    .A2(n_5228_o_0),
    .B(n_5092_o_0),
    .Y(n_5229_o_0));
 OAI31xp33_ASAP7_75t_R n_5230 (.A1(n_5216_o_0),
    .A2(n_5154_o_0),
    .A3(n_5159_o_0),
    .B(n_5009_o_0),
    .Y(n_5230_o_0));
 INVx1_ASAP7_75t_R n_5231 (.A(n_5230_o_0),
    .Y(n_5231_o_0));
 INVx1_ASAP7_75t_R n_5232 (.A(n_5033_o_0),
    .Y(n_5232_o_0));
 NAND3xp33_ASAP7_75t_R n_5233 (.A(n_5064_o_0),
    .B(n_5060_o_0),
    .C(n_5232_o_0),
    .Y(n_5233_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5234 (.A1(net60),
    .A2(n_4935_o_0),
    .B(n_5086_o_0),
    .C(n_5082_o_0),
    .Y(n_5234_o_0));
 OAI21xp33_ASAP7_75t_R n_5235 (.A1(n_4986_o_0),
    .A2(n_5234_o_0),
    .B(n_5092_o_0),
    .Y(n_5235_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5236 (.A1(n_5231_o_0),
    .A2(n_5233_o_0),
    .B(n_5235_o_0),
    .C(n_4832_o_0),
    .Y(n_5236_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5237 (.A1(n_5225_o_0),
    .A2(n_5226_o_0),
    .B(n_5229_o_0),
    .C(n_5236_o_0),
    .Y(n_5237_o_0));
 AOI31xp33_ASAP7_75t_R n_5238 (.A1(n_5084_o_0),
    .A2(n_5220_o_0),
    .A3(n_5224_o_0),
    .B(n_5237_o_0),
    .Y(n_5238_o_0));
 OAI21xp33_ASAP7_75t_R n_5239 (.A1(n_5167_o_0),
    .A2(n_5141_o_0),
    .B(n_5009_o_0),
    .Y(n_5239_o_0));
 AOI21xp33_ASAP7_75t_R n_5240 (.A1(n_4991_o_0),
    .A2(n_5087_o_0),
    .B(n_5239_o_0),
    .Y(n_5240_o_0));
 INVx1_ASAP7_75t_R n_5241 (.A(n_5115_o_0),
    .Y(n_5241_o_0));
 OAI21xp33_ASAP7_75t_R n_5242 (.A1(n_5062_o_0),
    .A2(n_5052_o_0),
    .B(n_5053_o_0),
    .Y(n_5242_o_0));
 AOI21xp33_ASAP7_75t_R n_5243 (.A1(n_5241_o_0),
    .A2(n_5022_o_0),
    .B(n_5242_o_0),
    .Y(n_5243_o_0));
 AOI22xp33_ASAP7_75t_R n_5244 (.A1(n_5027_o_0),
    .A2(n_5022_o_0),
    .B1(n_4858_o_0),
    .B2(n_5045_o_0),
    .Y(n_5244_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5245 (.A1(n_4859_o_0),
    .A2(n_4936_o_0),
    .B(n_5209_o_0),
    .C(n_5093_o_0),
    .Y(n_5245_o_0));
 OA21x2_ASAP7_75t_R n_5246 (.A1(n_4986_o_0),
    .A2(n_5244_o_0),
    .B(n_5245_o_0),
    .Y(n_5246_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5247 (.A1(n_5240_o_0),
    .A2(n_5243_o_0),
    .B(n_5093_o_0),
    .C(n_5246_o_0),
    .Y(n_5247_o_0));
 AOI21xp33_ASAP7_75t_R n_5248 (.A1(net60),
    .A2(n_4935_o_0),
    .B(n_5167_o_0),
    .Y(n_5248_o_0));
 AOI31xp33_ASAP7_75t_R n_5249 (.A1(n_4990_o_0),
    .A2(n_5051_o_0),
    .A3(n_4859_o_0),
    .B(n_5248_o_0),
    .Y(n_5249_o_0));
 INVx1_ASAP7_75t_R n_5250 (.A(n_5249_o_0),
    .Y(n_5250_o_0));
 AOI211xp5_ASAP7_75t_R n_5251 (.A1(n_5250_o_0),
    .A2(n_5009_o_0),
    .B(n_4811_o_0),
    .C(n_5205_o_0),
    .Y(n_5251_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5252 (.A1(n_4997_o_0),
    .A2(n_5001_o_0),
    .B(net95),
    .C(n_5114_o_0),
    .Y(n_5252_o_0));
 OAI21xp33_ASAP7_75t_R n_5253 (.A1(n_5070_o_0),
    .A2(n_4936_o_0),
    .B(n_4955_o_0),
    .Y(n_5253_o_0));
 OAI211xp5_ASAP7_75t_R n_5254 (.A1(n_5141_o_0),
    .A2(n_5086_o_0),
    .B(n_5253_o_0),
    .C(n_4970_o_0),
    .Y(n_5254_o_0));
 OAI32xp33_ASAP7_75t_R n_5255 (.A1(n_4810_o_0),
    .A2(n_4970_o_0),
    .A3(n_5252_o_0),
    .B1(n_5254_o_0),
    .B2(n_5093_o_0),
    .Y(n_5255_o_0));
 NOR3xp33_ASAP7_75t_R n_5256 (.A(n_5251_o_0),
    .B(n_5255_o_0),
    .C(n_5084_o_0),
    .Y(n_5256_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5257 (.A1(n_5015_o_0),
    .A2(n_5247_o_0),
    .B(n_5256_o_0),
    .C(n_4821_o_0),
    .Y(n_5257_o_0));
 OAI21xp33_ASAP7_75t_R n_5258 (.A1(n_4821_o_0),
    .A2(n_5238_o_0),
    .B(n_5257_o_0),
    .Y(n_5258_o_0));
 AOI21xp33_ASAP7_75t_R n_5259 (.A1(n_4998_o_0),
    .A2(net57),
    .B(n_4955_o_0),
    .Y(n_5259_o_0));
 AOI21xp33_ASAP7_75t_R n_5260 (.A1(n_5125_o_0),
    .A2(n_5259_o_0),
    .B(n_4986_o_0),
    .Y(n_5260_o_0));
 OAI31xp33_ASAP7_75t_R n_5261 (.A1(n_4859_o_0),
    .A2(n_5004_o_0),
    .A3(n_5033_o_0),
    .B(n_5260_o_0),
    .Y(n_5261_o_0));
 INVx1_ASAP7_75t_R n_5262 (.A(n_5261_o_0),
    .Y(n_5262_o_0));
 AOI211xp5_ASAP7_75t_R n_5263 (.A1(n_5017_o_0),
    .A2(n_5208_o_0),
    .B(n_5162_o_0),
    .C(n_4970_o_0),
    .Y(n_5263_o_0));
 AOI21xp33_ASAP7_75t_R n_5264 (.A1(n_5017_o_0),
    .A2(n_5001_o_0),
    .B(net95),
    .Y(n_5264_o_0));
 INVx1_ASAP7_75t_R n_5265 (.A(n_5046_o_0),
    .Y(n_5265_o_0));
 OAI211xp5_ASAP7_75t_R n_5266 (.A1(n_4998_o_0),
    .A2(net69),
    .B(n_5265_o_0),
    .C(n_4858_o_0),
    .Y(n_5266_o_0));
 OAI31xp33_ASAP7_75t_R n_5267 (.A1(n_4955_o_0),
    .A2(n_5055_o_0),
    .A3(n_5141_o_0),
    .B(n_5266_o_0),
    .Y(n_5267_o_0));
 OAI221xp5_ASAP7_75t_R n_5268 (.A1(n_5264_o_0),
    .A2(n_4996_o_0),
    .B1(n_4986_o_0),
    .B2(n_5267_o_0),
    .C(n_5084_o_0),
    .Y(n_5268_o_0));
 OAI31xp33_ASAP7_75t_R n_5269 (.A1(n_5015_o_0),
    .A2(n_5262_o_0),
    .A3(n_5263_o_0),
    .B(n_5268_o_0),
    .Y(n_5269_o_0));
 AOI21xp33_ASAP7_75t_R n_5270 (.A1(n_4810_o_0),
    .A2(n_5269_o_0),
    .B(n_5041_o_0),
    .Y(n_5270_o_0));
 AOI211xp5_ASAP7_75t_R n_5271 (.A1(n_4955_o_0),
    .A2(n_5008_o_0),
    .B(n_4982_o_0),
    .C(n_4936_o_0),
    .Y(n_5271_o_0));
 NAND2xp33_ASAP7_75t_R n_5272 (.A(n_4954_o_0),
    .B(n_5034_o_0),
    .Y(n_5272_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5273 (.A1(net60),
    .A2(n_5022_o_0),
    .B(n_5272_o_0),
    .C(n_5009_o_0),
    .Y(n_5273_o_0));
 AOI31xp33_ASAP7_75t_R n_5274 (.A1(n_4858_o_0),
    .A2(n_5265_o_0),
    .A3(n_5047_o_0),
    .B(n_5273_o_0),
    .Y(n_5274_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5275 (.A1(n_4970_o_0),
    .A2(n_5271_o_0),
    .B(n_5274_o_0),
    .C(n_5015_o_0),
    .Y(n_5275_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5276 (.A1(n_4858_o_0),
    .A2(n_5017_o_0),
    .B(n_5123_o_0),
    .C(n_5060_o_0),
    .Y(n_5276_o_0));
 AO21x1_ASAP7_75t_R n_5277 (.A1(n_5047_o_0),
    .A2(n_4858_o_0),
    .B(n_5045_o_0),
    .Y(n_5277_o_0));
 AOI21xp33_ASAP7_75t_R n_5278 (.A1(n_4970_o_0),
    .A2(n_5277_o_0),
    .B(n_5084_o_0),
    .Y(n_5278_o_0));
 OAI21xp33_ASAP7_75t_R n_5279 (.A1(net51),
    .A2(n_5276_o_0),
    .B(n_5278_o_0),
    .Y(n_5279_o_0));
 NAND3xp33_ASAP7_75t_R n_5280 (.A(n_5275_o_0),
    .B(n_5279_o_0),
    .C(n_5092_o_0),
    .Y(n_5280_o_0));
 NOR2xp33_ASAP7_75t_R n_5281 (.A(n_5026_o_0),
    .B(n_5116_o_0),
    .Y(n_5281_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5282 (.A1(n_4858_o_0),
    .A2(n_5232_o_0),
    .B(n_5281_o_0),
    .C(n_5047_o_0),
    .Y(n_5282_o_0));
 NOR2xp33_ASAP7_75t_R n_5283 (.A(n_4934_o_0),
    .B(n_4976_o_0),
    .Y(n_5283_o_0));
 OAI22xp33_ASAP7_75t_R n_5284 (.A1(n_5008_o_0),
    .A2(n_4859_o_0),
    .B1(n_4955_o_0),
    .B2(n_5283_o_0),
    .Y(n_5284_o_0));
 AOI21xp33_ASAP7_75t_R n_5285 (.A1(n_4986_o_0),
    .A2(n_5284_o_0),
    .B(n_5014_o_0),
    .Y(n_5285_o_0));
 OAI21xp33_ASAP7_75t_R n_5286 (.A1(n_4859_o_0),
    .A2(n_5168_o_0),
    .B(n_5133_o_0),
    .Y(n_5286_o_0));
 OAI31xp33_ASAP7_75t_R n_5287 (.A1(n_4985_o_0),
    .A2(n_5190_o_0),
    .A3(n_5055_o_0),
    .B(n_4992_o_0),
    .Y(n_5287_o_0));
 AOI211xp5_ASAP7_75t_R n_5288 (.A1(n_4970_o_0),
    .A2(n_5286_o_0),
    .B(n_5287_o_0),
    .C(n_5084_o_0),
    .Y(n_5288_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5289 (.A1(n_5009_o_0),
    .A2(n_5282_o_0),
    .B(n_5285_o_0),
    .C(n_5288_o_0),
    .Y(n_5289_o_0));
 AOI21xp33_ASAP7_75t_R n_5290 (.A1(n_5001_o_0),
    .A2(n_5123_o_0),
    .B(n_5083_o_0),
    .Y(n_5290_o_0));
 AOI21xp33_ASAP7_75t_R n_5291 (.A1(n_5061_o_0),
    .A2(n_5260_o_0),
    .B(n_4832_o_0),
    .Y(n_5291_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5292 (.A1(n_5001_o_0),
    .A2(n_5182_o_0),
    .B(n_4955_o_0),
    .C(n_5098_o_0),
    .Y(n_5292_o_0));
 AOI21xp33_ASAP7_75t_R n_5293 (.A1(n_4976_o_0),
    .A2(n_4954_o_0),
    .B(net60),
    .Y(n_5293_o_0));
 OAI21xp33_ASAP7_75t_R n_5294 (.A1(n_4858_o_0),
    .A2(n_5074_o_0),
    .B(n_4986_o_0),
    .Y(n_5294_o_0));
 OAI21xp33_ASAP7_75t_R n_5295 (.A1(n_5293_o_0),
    .A2(n_5294_o_0),
    .B(n_4832_o_0),
    .Y(n_5295_o_0));
 AOI21xp33_ASAP7_75t_R n_5296 (.A1(n_4970_o_0),
    .A2(n_5292_o_0),
    .B(n_5295_o_0),
    .Y(n_5296_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5297 (.A1(net51),
    .A2(n_5290_o_0),
    .B(n_5291_o_0),
    .C(n_5296_o_0),
    .Y(n_5297_o_0));
 AOI22xp33_ASAP7_75t_R n_5298 (.A1(n_5289_o_0),
    .A2(n_5092_o_0),
    .B1(n_4810_o_0),
    .B2(n_5297_o_0),
    .Y(n_5298_o_0));
 AOI22xp33_ASAP7_75t_R n_5299 (.A1(n_5270_o_0),
    .A2(n_5280_o_0),
    .B1(n_4821_o_0),
    .B2(n_5298_o_0),
    .Y(n_5299_o_0));
 AOI21xp33_ASAP7_75t_R n_5300 (.A1(n_4990_o_0),
    .A2(n_5105_o_0),
    .B(n_4982_o_0),
    .Y(n_5300_o_0));
 OAI21xp33_ASAP7_75t_R n_5301 (.A1(n_4976_o_0),
    .A2(n_5026_o_0),
    .B(n_5300_o_0),
    .Y(n_5301_o_0));
 INVx1_ASAP7_75t_R n_5302 (.A(n_5080_o_0),
    .Y(n_5302_o_0));
 NAND2xp33_ASAP7_75t_R n_5303 (.A(n_4899_o_0),
    .B(n_4858_o_0),
    .Y(n_5303_o_0));
 AOI211xp5_ASAP7_75t_R n_5304 (.A1(n_5302_o_0),
    .A2(n_5303_o_0),
    .B(n_5093_o_0),
    .C(n_4985_o_0),
    .Y(n_5304_o_0));
 AOI31xp33_ASAP7_75t_R n_5305 (.A1(n_4810_o_0),
    .A2(n_5301_o_0),
    .A3(n_4986_o_0),
    .B(n_5304_o_0),
    .Y(n_5305_o_0));
 AOI21xp33_ASAP7_75t_R n_5306 (.A1(n_5047_o_0),
    .A2(n_5259_o_0),
    .B(n_4810_o_0),
    .Y(n_5306_o_0));
 OAI21xp33_ASAP7_75t_R n_5307 (.A1(n_4956_o_0),
    .A2(n_5036_o_0),
    .B(n_5306_o_0),
    .Y(n_5307_o_0));
 AOI31xp33_ASAP7_75t_R n_5308 (.A1(n_4954_o_0),
    .A2(n_4990_o_0),
    .A3(n_5074_o_0),
    .B(n_5092_o_0),
    .Y(n_5308_o_0));
 OAI21xp33_ASAP7_75t_R n_5309 (.A1(n_5115_o_0),
    .A2(n_5029_o_0),
    .B(n_5308_o_0),
    .Y(n_5309_o_0));
 NAND3xp33_ASAP7_75t_R n_5310 (.A(n_5307_o_0),
    .B(n_5309_o_0),
    .C(n_4970_o_0),
    .Y(n_5310_o_0));
 OAI21xp33_ASAP7_75t_R n_5311 (.A1(n_4858_o_0),
    .A2(n_4981_o_0),
    .B(n_5075_o_0),
    .Y(n_5311_o_0));
 AOI311xp33_ASAP7_75t_R n_5312 (.A1(n_4954_o_0),
    .A2(n_5020_o_0),
    .A3(n_5074_o_0),
    .B(n_4811_o_0),
    .C(n_5009_o_0),
    .Y(n_5312_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5313 (.A1(n_4980_o_0),
    .A2(n_5029_o_0),
    .B(n_4956_o_0),
    .C(n_5312_o_0),
    .Y(n_5313_o_0));
 AOI22xp33_ASAP7_75t_R n_5314 (.A1(n_4990_o_0),
    .A2(n_4954_o_0),
    .B1(n_4858_o_0),
    .B2(n_4935_o_0),
    .Y(n_5314_o_0));
 NAND2xp33_ASAP7_75t_R n_5315 (.A(n_4954_o_0),
    .B(n_4990_o_0),
    .Y(n_5315_o_0));
 OAI21xp33_ASAP7_75t_R n_5316 (.A1(n_4872_o_0),
    .A2(n_5019_o_0),
    .B(n_4899_o_0),
    .Y(n_5316_o_0));
 AOI31xp33_ASAP7_75t_R n_5317 (.A1(n_4858_o_0),
    .A2(n_5092_o_0),
    .A3(n_5316_o_0),
    .B(n_4970_o_0),
    .Y(n_5317_o_0));
 OA21x2_ASAP7_75t_R n_5318 (.A1(n_5315_o_0),
    .A2(n_5036_o_0),
    .B(n_5317_o_0),
    .Y(n_5318_o_0));
 OAI21xp33_ASAP7_75t_R n_5319 (.A1(n_4811_o_0),
    .A2(n_5314_o_0),
    .B(n_5318_o_0),
    .Y(n_5319_o_0));
 OAI311xp33_ASAP7_75t_R n_5320 (.A1(n_4810_o_0),
    .A2(n_4986_o_0),
    .A3(n_5311_o_0),
    .B1(n_5313_o_0),
    .C1(n_5319_o_0),
    .Y(n_5320_o_0));
 AOI32xp33_ASAP7_75t_R n_5321 (.A1(n_4832_o_0),
    .A2(n_5305_o_0),
    .A3(n_5310_o_0),
    .B1(n_5320_o_0),
    .B2(n_5015_o_0),
    .Y(n_5321_o_0));
 AOI22xp33_ASAP7_75t_R n_5322 (.A1(n_5241_o_0),
    .A2(n_5081_o_0),
    .B1(n_5056_o_0),
    .B2(net95),
    .Y(n_5322_o_0));
 AO31x2_ASAP7_75t_R n_5323 (.A1(n_5253_o_0),
    .A2(n_5086_o_0),
    .A3(n_5009_o_0),
    .B(n_5092_o_0),
    .Y(n_5323_o_0));
 AOI21xp33_ASAP7_75t_R n_5324 (.A1(n_4970_o_0),
    .A2(n_5322_o_0),
    .B(n_5323_o_0),
    .Y(n_5324_o_0));
 AOI21xp33_ASAP7_75t_R n_5325 (.A1(n_4935_o_0),
    .A2(net60),
    .B(n_5046_o_0),
    .Y(n_5325_o_0));
 NOR3xp33_ASAP7_75t_R n_5326 (.A(n_5200_o_0),
    .B(n_4899_o_0),
    .C(n_4859_o_0),
    .Y(n_5326_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5327 (.A1(n_5325_o_0),
    .A2(net95),
    .B(n_5326_o_0),
    .C(n_4970_o_0),
    .Y(n_5327_o_0));
 AOI21xp33_ASAP7_75t_R n_5328 (.A1(n_5038_o_0),
    .A2(n_5327_o_0),
    .B(n_5093_o_0),
    .Y(n_5328_o_0));
 NAND3xp33_ASAP7_75t_R n_5329 (.A(n_4986_o_0),
    .B(n_5074_o_0),
    .C(n_4858_o_0),
    .Y(n_5329_o_0));
 OAI31xp33_ASAP7_75t_R n_5330 (.A1(n_5055_o_0),
    .A2(n_5329_o_0),
    .A3(n_5093_o_0),
    .B(n_4832_o_0),
    .Y(n_5330_o_0));
 NOR2xp33_ASAP7_75t_R n_5331 (.A(n_2521_o_0),
    .B(n_4965_o_0),
    .Y(n_5331_o_0));
 OAI321xp33_ASAP7_75t_R n_5332 (.A1(n_4999_o_0),
    .A2(n_4976_o_0),
    .A3(n_4974_o_0),
    .B1(n_4975_o_0),
    .B2(n_4952_o_0),
    .C(n_4954_o_0),
    .Y(n_5332_o_0));
 OAI31xp33_ASAP7_75t_R n_5333 (.A1(n_4999_o_0),
    .A2(n_4974_o_0),
    .A3(n_4859_o_0),
    .B(n_5332_o_0),
    .Y(n_5333_o_0));
 OA21x2_ASAP7_75t_R n_5334 (.A1(n_4984_o_0),
    .A2(n_5331_o_0),
    .B(n_5333_o_0),
    .Y(n_5334_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5335 (.A1(n_4990_o_0),
    .A2(n_5051_o_0),
    .B(n_4859_o_0),
    .C(n_4985_o_0),
    .Y(n_5335_o_0));
 AOI21xp33_ASAP7_75t_R n_5336 (.A1(n_5071_o_0),
    .A2(n_5125_o_0),
    .B(n_5335_o_0),
    .Y(n_5336_o_0));
 NOR3xp33_ASAP7_75t_R n_5337 (.A(net57),
    .B(n_4898_o_0),
    .C(n_4949_o_0),
    .Y(n_5337_o_0));
 NOR5xp2_ASAP7_75t_R n_5338 (.A(n_5337_o_0),
    .B(n_5003_o_0),
    .C(n_4954_o_0),
    .D(n_4985_o_0),
    .E(n_5007_o_0),
    .Y(n_5338_o_0));
 AOI211xp5_ASAP7_75t_R n_5339 (.A1(n_5000_o_0),
    .A2(net60),
    .B(n_5062_o_0),
    .C(n_4858_o_0),
    .Y(n_5339_o_0));
 AOI22xp33_ASAP7_75t_R n_5340 (.A1(n_5008_o_0),
    .A2(n_4955_o_0),
    .B1(n_5339_o_0),
    .B2(n_4985_o_0),
    .Y(n_5340_o_0));
 OAI21xp33_ASAP7_75t_R n_5341 (.A1(n_5157_o_0),
    .A2(n_4956_o_0),
    .B(n_5197_o_0),
    .Y(n_5341_o_0));
 OAI221xp5_ASAP7_75t_R n_5342 (.A1(n_5338_o_0),
    .A2(n_5340_o_0),
    .B1(n_4970_o_0),
    .B2(n_5341_o_0),
    .C(n_4810_o_0),
    .Y(n_5342_o_0));
 OAI31xp33_ASAP7_75t_R n_5343 (.A1(n_5093_o_0),
    .A2(n_5334_o_0),
    .A3(n_5336_o_0),
    .B(n_5342_o_0),
    .Y(n_5343_o_0));
 OAI21xp33_ASAP7_75t_R n_5344 (.A1(n_4831_o_0),
    .A2(n_4829_o_0),
    .B(n_5343_o_0),
    .Y(n_5344_o_0));
 OAI31xp33_ASAP7_75t_R n_5345 (.A1(n_5324_o_0),
    .A2(n_5328_o_0),
    .A3(n_5330_o_0),
    .B(n_5344_o_0),
    .Y(n_5345_o_0));
 OAI21xp33_ASAP7_75t_R n_5346 (.A1(n_4818_o_0),
    .A2(n_4820_o_0),
    .B(n_5345_o_0),
    .Y(n_5346_o_0));
 OA21x2_ASAP7_75t_R n_5347 (.A1(n_4822_o_0),
    .A2(n_5321_o_0),
    .B(n_5346_o_0),
    .Y(n_5347_o_0));
 AND3x1_ASAP7_75t_R n_5348 (.A(n_5189_o_0),
    .B(n_5316_o_0),
    .C(net95),
    .Y(n_5348_o_0));
 AOI31xp33_ASAP7_75t_R n_5349 (.A1(n_4858_o_0),
    .A2(n_4997_o_0),
    .A3(n_5265_o_0),
    .B(n_5348_o_0),
    .Y(n_5349_o_0));
 NAND3xp33_ASAP7_75t_R n_5350 (.A(n_5158_o_0),
    .B(n_5020_o_0),
    .C(net95),
    .Y(n_5350_o_0));
 OAI31xp33_ASAP7_75t_R n_5351 (.A1(n_4859_o_0),
    .A2(n_5036_o_0),
    .A3(n_5033_o_0),
    .B(n_5350_o_0),
    .Y(n_5351_o_0));
 AOI21xp33_ASAP7_75t_R n_5352 (.A1(n_5092_o_0),
    .A2(n_5351_o_0),
    .B(n_4970_o_0),
    .Y(n_5352_o_0));
 OAI21xp33_ASAP7_75t_R n_5353 (.A1(n_4811_o_0),
    .A2(n_5349_o_0),
    .B(n_5352_o_0),
    .Y(n_5353_o_0));
 NAND3xp33_ASAP7_75t_R n_5354 (.A(n_5017_o_0),
    .B(n_5081_o_0),
    .C(n_4858_o_0),
    .Y(n_5354_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5355 (.A1(n_5029_o_0),
    .A2(n_5028_o_0),
    .B(n_5354_o_0),
    .C(n_4811_o_0),
    .Y(n_5355_o_0));
 INVx1_ASAP7_75t_R n_5356 (.A(n_5355_o_0),
    .Y(n_5356_o_0));
 NAND2xp33_ASAP7_75t_R n_5357 (.A(n_4998_o_0),
    .B(n_5022_o_0),
    .Y(n_5357_o_0));
 OAI211xp5_ASAP7_75t_R n_5358 (.A1(n_4858_o_0),
    .A2(n_5357_o_0),
    .B(n_5174_o_0),
    .C(n_5092_o_0),
    .Y(n_5358_o_0));
 NAND3xp33_ASAP7_75t_R n_5359 (.A(n_5356_o_0),
    .B(n_5358_o_0),
    .C(net51),
    .Y(n_5359_o_0));
 NAND3xp33_ASAP7_75t_R n_5360 (.A(n_5047_o_0),
    .B(n_5034_o_0),
    .C(net95),
    .Y(n_5360_o_0));
 OAI31xp33_ASAP7_75t_R n_5361 (.A1(n_4859_o_0),
    .A2(n_5057_o_0),
    .A3(n_5168_o_0),
    .B(n_5360_o_0),
    .Y(n_5361_o_0));
 AOI211xp5_ASAP7_75t_R n_5362 (.A1(n_4976_o_0),
    .A2(net60),
    .B(n_4936_o_0),
    .C(n_4859_o_0),
    .Y(n_5362_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5363 (.A1(n_5189_o_0),
    .A2(n_5196_o_0),
    .B(n_4858_o_0),
    .C(n_4970_o_0),
    .Y(n_5363_o_0));
 OAI21xp33_ASAP7_75t_R n_5364 (.A1(n_5362_o_0),
    .A2(n_5363_o_0),
    .B(n_5093_o_0),
    .Y(n_5364_o_0));
 AOI21xp33_ASAP7_75t_R n_5365 (.A1(n_4986_o_0),
    .A2(n_5361_o_0),
    .B(n_5364_o_0),
    .Y(n_5365_o_0));
 OAI21xp33_ASAP7_75t_R n_5366 (.A1(n_5004_o_0),
    .A2(n_4936_o_0),
    .B(n_4955_o_0),
    .Y(n_5366_o_0));
 OAI21xp33_ASAP7_75t_R n_5367 (.A1(n_4858_o_0),
    .A2(n_5001_o_0),
    .B(n_5366_o_0),
    .Y(n_5367_o_0));
 NAND2xp33_ASAP7_75t_R n_5368 (.A(net57),
    .B(n_4859_o_0),
    .Y(n_5368_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5369 (.A1(n_5154_o_0),
    .A2(n_5116_o_0),
    .B(n_5368_o_0),
    .C(n_4970_o_0),
    .Y(n_5369_o_0));
 AOI211xp5_ASAP7_75t_R n_5370 (.A1(n_5367_o_0),
    .A2(net51),
    .B(n_5093_o_0),
    .C(n_5369_o_0),
    .Y(n_5370_o_0));
 NOR3xp33_ASAP7_75t_R n_5371 (.A(n_5365_o_0),
    .B(n_5370_o_0),
    .C(n_5015_o_0),
    .Y(n_5371_o_0));
 AOI31xp33_ASAP7_75t_R n_5372 (.A1(n_5084_o_0),
    .A2(n_5353_o_0),
    .A3(n_5359_o_0),
    .B(n_5371_o_0),
    .Y(n_5372_o_0));
 AND2x2_ASAP7_75t_R n_5373 (.A(n_4986_o_0),
    .B(n_5192_o_0),
    .Y(n_5373_o_0));
 NOR2xp33_ASAP7_75t_R n_5374 (.A(n_4811_o_0),
    .B(n_5009_o_0),
    .Y(n_5374_o_0));
 OA211x2_ASAP7_75t_R n_5375 (.A1(n_5033_o_0),
    .A2(n_5048_o_0),
    .B(n_5374_o_0),
    .C(n_5052_o_0),
    .Y(n_5375_o_0));
 AOI31xp33_ASAP7_75t_R n_5376 (.A1(n_4858_o_0),
    .A2(n_5020_o_0),
    .A3(n_5074_o_0),
    .B(n_4986_o_0),
    .Y(n_5376_o_0));
 OAI21xp33_ASAP7_75t_R n_5377 (.A1(n_5129_o_0),
    .A2(n_4955_o_0),
    .B(n_5376_o_0),
    .Y(n_5377_o_0));
 XNOR2xp5_ASAP7_75t_R n_5378 (.A(net57),
    .B(net60),
    .Y(n_5378_o_0));
 AOI21xp33_ASAP7_75t_R n_5379 (.A1(n_5047_o_0),
    .A2(n_5259_o_0),
    .B(n_4970_o_0),
    .Y(n_5379_o_0));
 OAI21xp33_ASAP7_75t_R n_5380 (.A1(n_4859_o_0),
    .A2(n_5378_o_0),
    .B(n_5379_o_0),
    .Y(n_5380_o_0));
 AOI21xp33_ASAP7_75t_R n_5381 (.A1(n_5377_o_0),
    .A2(n_5380_o_0),
    .B(n_4810_o_0),
    .Y(n_5381_o_0));
 AOI211xp5_ASAP7_75t_R n_5382 (.A1(n_4810_o_0),
    .A2(n_5373_o_0),
    .B(n_5375_o_0),
    .C(n_5381_o_0),
    .Y(n_5382_o_0));
 OAI21xp33_ASAP7_75t_R n_5383 (.A1(net60),
    .A2(n_5283_o_0),
    .B(n_4859_o_0),
    .Y(n_5383_o_0));
 OAI211xp5_ASAP7_75t_R n_5384 (.A1(net57),
    .A2(net95),
    .B(n_5383_o_0),
    .C(n_5303_o_0),
    .Y(n_5384_o_0));
 INVx1_ASAP7_75t_R n_5385 (.A(n_5303_o_0),
    .Y(n_5385_o_0));
 OAI211xp5_ASAP7_75t_R n_5386 (.A1(n_5385_o_0),
    .A2(net69),
    .B(n_4986_o_0),
    .C(n_4997_o_0),
    .Y(n_5386_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5387 (.A1(n_5384_o_0),
    .A2(n_5129_o_0),
    .B(n_5009_o_0),
    .C(n_5386_o_0),
    .Y(n_5387_o_0));
 AOI21xp33_ASAP7_75t_R n_5388 (.A1(n_4954_o_0),
    .A2(n_5020_o_0),
    .B(n_4970_o_0),
    .Y(n_5388_o_0));
 OAI311xp33_ASAP7_75t_R n_5389 (.A1(n_4859_o_0),
    .A2(n_5070_o_0),
    .A3(n_4936_o_0),
    .B1(n_5093_o_0),
    .C1(n_5388_o_0),
    .Y(n_5389_o_0));
 OA21x2_ASAP7_75t_R n_5390 (.A1(n_5387_o_0),
    .A2(n_4810_o_0),
    .B(n_5389_o_0),
    .Y(n_5390_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5391 (.A1(n_5060_o_0),
    .A2(n_5073_o_0),
    .B(n_5144_o_0),
    .C(n_5374_o_0),
    .Y(n_5391_o_0));
 AOI31xp33_ASAP7_75t_R n_5392 (.A1(n_5014_o_0),
    .A2(n_5390_o_0),
    .A3(n_5391_o_0),
    .B(n_4822_o_0),
    .Y(n_5392_o_0));
 OAI21xp33_ASAP7_75t_R n_5393 (.A1(n_4832_o_0),
    .A2(n_5382_o_0),
    .B(n_5392_o_0),
    .Y(n_5393_o_0));
 OAI21xp33_ASAP7_75t_R n_5394 (.A1(n_4821_o_0),
    .A2(n_5372_o_0),
    .B(n_5393_o_0),
    .Y(n_5394_o_0));
 OAI21xp33_ASAP7_75t_R n_5395 (.A1(n_5059_o_0),
    .A2(n_5154_o_0),
    .B(n_5093_o_0),
    .Y(n_5395_o_0));
 AOI31xp33_ASAP7_75t_R n_5396 (.A1(net95),
    .A2(n_5034_o_0),
    .A3(n_5047_o_0),
    .B(n_5395_o_0),
    .Y(n_5396_o_0));
 OAI21xp33_ASAP7_75t_R n_5397 (.A1(n_5033_o_0),
    .A2(n_5048_o_0),
    .B(n_4811_o_0),
    .Y(n_5397_o_0));
 AOI21xp33_ASAP7_75t_R n_5398 (.A1(net95),
    .A2(n_5034_o_0),
    .B(n_5397_o_0),
    .Y(n_5398_o_0));
 OAI21xp33_ASAP7_75t_R n_5399 (.A1(n_5396_o_0),
    .A2(n_5398_o_0),
    .B(n_5009_o_0),
    .Y(n_5399_o_0));
 AOI21xp33_ASAP7_75t_R n_5400 (.A1(n_5034_o_0),
    .A2(n_5023_o_0),
    .B(n_5092_o_0),
    .Y(n_5400_o_0));
 OA21x2_ASAP7_75t_R n_5401 (.A1(n_5070_o_0),
    .A2(n_5086_o_0),
    .B(n_5400_o_0),
    .Y(n_5401_o_0));
 AOI21xp33_ASAP7_75t_R n_5402 (.A1(n_5071_o_0),
    .A2(n_5265_o_0),
    .B(n_4810_o_0),
    .Y(n_5402_o_0));
 OAI21xp33_ASAP7_75t_R n_5403 (.A1(n_5115_o_0),
    .A2(n_4899_o_0),
    .B(n_5402_o_0),
    .Y(n_5403_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5404 (.A1(n_5057_o_0),
    .A2(n_5203_o_0),
    .B(n_4858_o_0),
    .C(n_5403_o_0),
    .Y(n_5404_o_0));
 OAI21xp33_ASAP7_75t_R n_5405 (.A1(n_5401_o_0),
    .A2(n_5404_o_0),
    .B(net51),
    .Y(n_5405_o_0));
 AOI21xp33_ASAP7_75t_R n_5406 (.A1(n_5399_o_0),
    .A2(n_5405_o_0),
    .B(n_4822_o_0),
    .Y(n_5406_o_0));
 OAI211xp5_ASAP7_75t_R n_5407 (.A1(net95),
    .A2(n_5182_o_0),
    .B(n_5005_o_0),
    .C(n_5001_o_0),
    .Y(n_5407_o_0));
 NOR3xp33_ASAP7_75t_R n_5408 (.A(n_5057_o_0),
    .B(n_5070_o_0),
    .C(n_5203_o_0),
    .Y(n_5408_o_0));
 AOI31xp33_ASAP7_75t_R n_5409 (.A1(n_4858_o_0),
    .A2(n_5020_o_0),
    .A3(n_5051_o_0),
    .B(n_5093_o_0),
    .Y(n_5409_o_0));
 OAI21xp33_ASAP7_75t_R n_5410 (.A1(n_4858_o_0),
    .A2(n_5408_o_0),
    .B(n_5409_o_0),
    .Y(n_5410_o_0));
 OA21x2_ASAP7_75t_R n_5411 (.A1(n_4811_o_0),
    .A2(n_5407_o_0),
    .B(n_5410_o_0),
    .Y(n_5411_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5412 (.A1(n_4998_o_0),
    .A2(n_4899_o_0),
    .B(net69),
    .C(n_4955_o_0),
    .Y(n_5412_o_0));
 OAI221xp5_ASAP7_75t_R n_5413 (.A1(n_4858_o_0),
    .A2(n_4993_o_0),
    .B1(n_5116_o_0),
    .B2(n_5154_o_0),
    .C(n_5093_o_0),
    .Y(n_5413_o_0));
 OAI31xp33_ASAP7_75t_R n_5414 (.A1(n_5093_o_0),
    .A2(n_5248_o_0),
    .A3(n_5412_o_0),
    .B(n_5413_o_0),
    .Y(n_5414_o_0));
 OAI21xp33_ASAP7_75t_R n_5415 (.A1(n_4986_o_0),
    .A2(n_5414_o_0),
    .B(n_4822_o_0),
    .Y(n_5415_o_0));
 AOI21xp33_ASAP7_75t_R n_5416 (.A1(n_5009_o_0),
    .A2(n_5411_o_0),
    .B(n_5415_o_0),
    .Y(n_5416_o_0));
 NAND2xp33_ASAP7_75t_R n_5417 (.A(n_5020_o_0),
    .B(n_5023_o_0),
    .Y(n_5417_o_0));
 OAI31xp33_ASAP7_75t_R n_5418 (.A1(n_4955_o_0),
    .A2(n_5070_o_0),
    .A3(n_5033_o_0),
    .B(n_5417_o_0),
    .Y(n_5418_o_0));
 NAND2xp33_ASAP7_75t_R n_5419 (.A(n_4810_o_0),
    .B(n_5418_o_0),
    .Y(n_5419_o_0));
 OAI31xp33_ASAP7_75t_R n_5420 (.A1(n_4955_o_0),
    .A2(n_5018_o_0),
    .A3(n_5116_o_0),
    .B(n_5098_o_0),
    .Y(n_5420_o_0));
 NAND2xp33_ASAP7_75t_R n_5421 (.A(n_5092_o_0),
    .B(n_5420_o_0),
    .Y(n_5421_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5422 (.A1(n_5022_o_0),
    .A2(net60),
    .B(n_4936_o_0),
    .C(n_4859_o_0),
    .Y(n_5422_o_0));
 OAI21xp33_ASAP7_75t_R n_5423 (.A1(net95),
    .A2(n_5101_o_0),
    .B(n_5422_o_0),
    .Y(n_5423_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5424 (.A1(n_4859_o_0),
    .A2(n_5283_o_0),
    .B(n_5005_o_0),
    .C(n_4810_o_0),
    .Y(n_5424_o_0));
 AOI211xp5_ASAP7_75t_R n_5425 (.A1(n_5423_o_0),
    .A2(n_5093_o_0),
    .B(n_4985_o_0),
    .C(n_5424_o_0),
    .Y(n_5425_o_0));
 AOI31xp33_ASAP7_75t_R n_5426 (.A1(n_4970_o_0),
    .A2(n_5419_o_0),
    .A3(n_5421_o_0),
    .B(n_5425_o_0),
    .Y(n_5426_o_0));
 AOI21xp33_ASAP7_75t_R n_5427 (.A1(n_5022_o_0),
    .A2(n_5027_o_0),
    .B(n_5092_o_0),
    .Y(n_5427_o_0));
 AOI211xp5_ASAP7_75t_R n_5428 (.A1(n_5259_o_0),
    .A2(n_5085_o_0),
    .B(n_5162_o_0),
    .C(n_4810_o_0),
    .Y(n_5428_o_0));
 AOI21xp33_ASAP7_75t_R n_5429 (.A1(n_5126_o_0),
    .A2(n_5427_o_0),
    .B(n_5428_o_0),
    .Y(n_5429_o_0));
 AOI31xp33_ASAP7_75t_R n_5430 (.A1(n_4954_o_0),
    .A2(n_5020_o_0),
    .A3(n_5085_o_0),
    .B(n_5092_o_0),
    .Y(n_5430_o_0));
 OA21x2_ASAP7_75t_R n_5431 (.A1(n_4859_o_0),
    .A2(n_5046_o_0),
    .B(n_5430_o_0),
    .Y(n_5431_o_0));
 NAND3xp33_ASAP7_75t_R n_5432 (.A(n_5017_o_0),
    .B(n_5060_o_0),
    .C(n_4858_o_0),
    .Y(n_5432_o_0));
 AOI21xp33_ASAP7_75t_R n_5433 (.A1(net95),
    .A2(n_4976_o_0),
    .B(n_4986_o_0),
    .Y(n_5433_o_0));
 AOI21xp33_ASAP7_75t_R n_5434 (.A1(n_5432_o_0),
    .A2(n_5433_o_0),
    .B(n_5374_o_0),
    .Y(n_5434_o_0));
 OAI21xp33_ASAP7_75t_R n_5435 (.A1(n_5431_o_0),
    .A2(n_5434_o_0),
    .B(n_4821_o_0),
    .Y(n_5435_o_0));
 AO21x1_ASAP7_75t_R n_5436 (.A1(n_4986_o_0),
    .A2(n_5429_o_0),
    .B(n_5435_o_0),
    .Y(n_5436_o_0));
 OAI211xp5_ASAP7_75t_R n_5437 (.A1(n_5426_o_0),
    .A2(n_4821_o_0),
    .B(n_5436_o_0),
    .C(n_5015_o_0),
    .Y(n_5437_o_0));
 OAI31xp33_ASAP7_75t_R n_5438 (.A1(n_5015_o_0),
    .A2(n_5406_o_0),
    .A3(n_5416_o_0),
    .B(n_5437_o_0),
    .Y(n_5438_o_0));
 XOR2xp5_ASAP7_75t_R n_5439 (.A(_01003_),
    .B(n_3012_o_0),
    .Y(n_5439_o_0));
 NOR2xp33_ASAP7_75t_R n_5440 (.A(n_3136_o_0),
    .B(n_5439_o_0),
    .Y(n_5440_o_0));
 NOR2xp33_ASAP7_75t_R n_5441 (.A(_00654_),
    .B(net),
    .Y(n_5441_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5442 (.A1(n_3136_o_0),
    .A2(n_5439_o_0),
    .B(n_5440_o_0),
    .C(net),
    .D(n_5441_o_0),
    .Y(n_5442_o_0));
 XNOR2xp5_ASAP7_75t_R n_5443 (.A(_00883_),
    .B(n_5442_o_0),
    .Y(n_5443_o_0));
 XNOR2xp5_ASAP7_75t_R n_5444 (.A(_00643_),
    .B(_01076_),
    .Y(n_5444_o_0));
 XOR2xp5_ASAP7_75t_R n_5445 (.A(_01077_),
    .B(_01116_),
    .Y(n_5445_o_0));
 XNOR2xp5_ASAP7_75t_R n_5446 (.A(n_5444_o_0),
    .B(n_5445_o_0),
    .Y(n_5446_o_0));
 XNOR2xp5_ASAP7_75t_R n_5447 (.A(_00997_),
    .B(n_3062_o_0),
    .Y(n_5447_o_0));
 XOR2xp5_ASAP7_75t_R n_5448 (.A(_00643_),
    .B(_01076_),
    .Y(n_5448_o_0));
 NAND2xp33_ASAP7_75t_R n_5449 (.A(n_5448_o_0),
    .B(n_5445_o_0),
    .Y(n_5449_o_0));
 XNOR2xp5_ASAP7_75t_R n_5450 (.A(_01077_),
    .B(_01116_),
    .Y(n_5450_o_0));
 NAND2xp33_ASAP7_75t_R n_5451 (.A(n_5444_o_0),
    .B(n_5450_o_0),
    .Y(n_5451_o_0));
 NAND2xp33_ASAP7_75t_R n_5452 (.A(_00997_),
    .B(n_3078_o_0),
    .Y(n_5452_o_0));
 INVx1_ASAP7_75t_R n_5453 (.A(_00997_),
    .Y(n_5453_o_0));
 NAND2xp33_ASAP7_75t_R n_5454 (.A(n_5453_o_0),
    .B(n_3062_o_0),
    .Y(n_5454_o_0));
 AOI22xp33_ASAP7_75t_R n_5455 (.A1(n_5449_o_0),
    .A2(n_5451_o_0),
    .B1(n_5452_o_0),
    .B2(n_5454_o_0),
    .Y(n_5455_o_0));
 NOR2xp33_ASAP7_75t_R n_5456 (.A(_00529_),
    .B(_00858_),
    .Y(n_5456_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5457 (.A1(n_5446_o_0),
    .A2(n_5447_o_0),
    .B(n_5455_o_0),
    .C(_00858_),
    .D(n_5456_o_0),
    .Y(n_5457_o_0));
 NAND2xp33_ASAP7_75t_R n_5458 (.A(_00877_),
    .B(n_5457_o_0),
    .Y(n_5458_o_0));
 OAI21x1_ASAP7_75t_R n_5459 (.A1(_00877_),
    .A2(n_5457_o_0),
    .B(n_5458_o_0),
    .Y(n_5459_o_0));
 INVx1_ASAP7_75t_R n_5460 (.A(_00998_),
    .Y(n_5460_o_0));
 NOR2xp33_ASAP7_75t_R n_5461 (.A(n_5460_o_0),
    .B(n_3037_o_0),
    .Y(n_5461_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5462 (.A1(n_3037_o_0),
    .A2(n_5460_o_0),
    .B(n_5461_o_0),
    .C(n_3080_o_0),
    .Y(n_5462_o_0));
 NAND2xp33_ASAP7_75t_R n_5463 (.A(n_5460_o_0),
    .B(n_3037_o_0),
    .Y(n_5463_o_0));
 OAI211xp5_ASAP7_75t_R n_5464 (.A1(n_3037_o_0),
    .A2(n_5460_o_0),
    .B(n_5463_o_0),
    .C(n_3063_o_0),
    .Y(n_5464_o_0));
 OR2x2_ASAP7_75t_R n_5465 (.A(_00532_),
    .B(_00858_),
    .Y(n_5465_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5466 (.A1(n_5462_o_0),
    .A2(n_5464_o_0),
    .B(n_3021_o_0),
    .C(n_5465_o_0),
    .Y(n_5466_o_0));
 NOR2xp33_ASAP7_75t_R n_5467 (.A(_00878_),
    .B(n_5466_o_0),
    .Y(n_5467_o_0));
 INVx1_ASAP7_75t_R n_5468 (.A(_00878_),
    .Y(n_5468_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5469 (.A1(n_5464_o_0),
    .A2(n_5462_o_0),
    .B(n_3021_o_0),
    .C(n_5465_o_0),
    .D(n_5468_o_0),
    .Y(n_5469_o_0));
 INVx1_ASAP7_75t_R n_5470 (.A(_00996_),
    .Y(n_5470_o_0));
 XOR2xp5_ASAP7_75t_R n_5471 (.A(_01043_),
    .B(_01115_),
    .Y(n_5471_o_0));
 NAND2xp33_ASAP7_75t_R n_5472 (.A(_01043_),
    .B(_01115_),
    .Y(n_5472_o_0));
 OAI211xp5_ASAP7_75t_R n_5473 (.A1(_01043_),
    .A2(_01115_),
    .B(n_5472_o_0),
    .C(n_5470_o_0),
    .Y(n_5473_o_0));
 OAI21xp33_ASAP7_75t_R n_5474 (.A1(n_5470_o_0),
    .A2(n_5471_o_0),
    .B(n_5473_o_0),
    .Y(n_5474_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5475 (.A1(_01043_),
    .A2(_01115_),
    .B(n_5472_o_0),
    .C(n_5470_o_0),
    .Y(n_5475_o_0));
 AOI211xp5_ASAP7_75t_R n_5476 (.A1(n_5471_o_0),
    .A2(n_5470_o_0),
    .B(n_5448_o_0),
    .C(n_5475_o_0),
    .Y(n_5476_o_0));
 NOR2xp33_ASAP7_75t_R n_5477 (.A(_00530_),
    .B(_00858_),
    .Y(n_5477_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5478 (.A1(n_5448_o_0),
    .A2(n_5474_o_0),
    .B(n_5476_o_0),
    .C(net39),
    .D(n_5477_o_0),
    .Y(n_5478_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5479 (.A1(n_5471_o_0),
    .A2(n_5470_o_0),
    .B(n_5475_o_0),
    .C(n_5448_o_0),
    .Y(n_5479_o_0));
 OAI211xp5_ASAP7_75t_R n_5480 (.A1(n_5471_o_0),
    .A2(n_5470_o_0),
    .B(n_5473_o_0),
    .C(n_5444_o_0),
    .Y(n_5480_o_0));
 INVx1_ASAP7_75t_R n_5481 (.A(n_5477_o_0),
    .Y(n_5481_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5482 (.A1(n_5479_o_0),
    .A2(n_5480_o_0),
    .B(net5),
    .C(n_5481_o_0),
    .D(_00876_),
    .Y(n_5482_o_0));
 AO21x1_ASAP7_75t_R n_5483 (.A1(_00876_),
    .A2(n_5478_o_0),
    .B(n_5482_o_0),
    .Y(n_5483_o_0));
 INVx2_ASAP7_75t_R n_5484 (.A(n_5483_o_0),
    .Y(n_5484_o_0));
 OAI21xp33_ASAP7_75t_R n_5485 (.A1(n_5467_o_0),
    .A2(n_5469_o_0),
    .B(n_5484_o_0),
    .Y(n_5485_o_0));
 NOR2xp33_ASAP7_75t_R n_5486 (.A(n_5459_o_0),
    .B(n_5485_o_0),
    .Y(n_5486_o_0));
 INVx1_ASAP7_75t_R n_5487 (.A(n_5486_o_0),
    .Y(n_5487_o_0));
 INVx1_ASAP7_75t_R n_5488 (.A(n_5466_o_0),
    .Y(n_5488_o_0));
 AOI21x1_ASAP7_75t_R n_5489 (.A1(n_5468_o_0),
    .A2(n_5488_o_0),
    .B(n_5469_o_0),
    .Y(n_5489_o_0));
 NAND2xp33_ASAP7_75t_R n_5490 (.A(n_5483_o_0),
    .B(n_5489_o_0),
    .Y(n_5490_o_0));
 XOR2xp5_ASAP7_75t_R n_5491 (.A(_00643_),
    .B(_01078_),
    .Y(n_5491_o_0));
 NAND2xp33_ASAP7_75t_R n_5492 (.A(n_3026_o_0),
    .B(n_5491_o_0),
    .Y(n_5492_o_0));
 OAI21xp33_ASAP7_75t_R n_5493 (.A1(n_3026_o_0),
    .A2(n_5491_o_0),
    .B(n_5492_o_0),
    .Y(n_5493_o_0));
 NAND2xp33_ASAP7_75t_R n_5494 (.A(_00999_),
    .B(n_3025_o_0),
    .Y(n_5494_o_0));
 OAI21xp33_ASAP7_75t_R n_5495 (.A1(_00999_),
    .A2(n_3025_o_0),
    .B(n_5494_o_0),
    .Y(n_5495_o_0));
 NAND2xp33_ASAP7_75t_R n_5496 (.A(n_5495_o_0),
    .B(n_5493_o_0),
    .Y(n_5496_o_0));
 OAI21xp33_ASAP7_75t_R n_5497 (.A1(n_5493_o_0),
    .A2(n_5495_o_0),
    .B(n_5496_o_0),
    .Y(n_5497_o_0));
 NOR2xp33_ASAP7_75t_R n_5498 (.A(_00658_),
    .B(_00858_),
    .Y(n_5498_o_0));
 AO21x1_ASAP7_75t_R n_5499 (.A1(n_5497_o_0),
    .A2(net),
    .B(n_5498_o_0),
    .Y(n_5499_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5500 (.A1(n_5497_o_0),
    .A2(net),
    .B(n_5498_o_0),
    .C(_00879_),
    .Y(n_5500_o_0));
 OAI21xp5_ASAP7_75t_R n_5501 (.A1(_00879_),
    .A2(n_5499_o_0),
    .B(n_5500_o_0),
    .Y(n_5501_o_0));
 NAND2xp33_ASAP7_75t_R n_5502 (.A(n_5490_o_0),
    .B(n_5501_o_0),
    .Y(n_5502_o_0));
 INVx1_ASAP7_75t_R n_5503 (.A(n_5502_o_0),
    .Y(n_5503_o_0));
 INVx1_ASAP7_75t_R n_5504 (.A(n_3005_o_0),
    .Y(n_5504_o_0));
 XNOR2xp5_ASAP7_75t_R n_5505 (.A(_01001_),
    .B(_01040_),
    .Y(n_5505_o_0));
 XNOR2xp5_ASAP7_75t_R n_5506 (.A(_01080_),
    .B(n_5505_o_0),
    .Y(n_5506_o_0));
 XNOR2xp5_ASAP7_75t_R n_5507 (.A(n_5504_o_0),
    .B(n_5506_o_0),
    .Y(n_5507_o_0));
 NOR2xp33_ASAP7_75t_R n_5508 (.A(_00656_),
    .B(net),
    .Y(n_5508_o_0));
 AOI21xp33_ASAP7_75t_R n_5509 (.A1(net39),
    .A2(n_5507_o_0),
    .B(n_5508_o_0),
    .Y(n_5509_o_0));
 XOR2xp5_ASAP7_75t_R n_5510 (.A(_00881_),
    .B(n_5509_o_0),
    .Y(n_5510_o_0));
 AOI21xp33_ASAP7_75t_R n_5511 (.A1(n_5487_o_0),
    .A2(n_5503_o_0),
    .B(n_5510_o_0),
    .Y(n_5511_o_0));
 INVx1_ASAP7_75t_R n_5512 (.A(_00879_),
    .Y(n_5512_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5513 (.A1(n_5497_o_0),
    .A2(net),
    .B(n_5498_o_0),
    .C(n_5512_o_0),
    .Y(n_5513_o_0));
 OAI21xp5_ASAP7_75t_R n_5514 (.A1(n_5512_o_0),
    .A2(n_5499_o_0),
    .B(n_5513_o_0),
    .Y(n_5514_o_0));
 OAI211xp5_ASAP7_75t_R n_5515 (.A1(n_5483_o_0),
    .A2(n_5489_o_0),
    .B(n_5514_o_0),
    .C(n_5459_o_0),
    .Y(n_5515_o_0));
 XNOR2xp5_ASAP7_75t_R n_5516 (.A(_00643_),
    .B(_01079_),
    .Y(n_5516_o_0));
 XOR2xp5_ASAP7_75t_R n_5517 (.A(n_3113_o_0),
    .B(n_5516_o_0),
    .Y(n_5517_o_0));
 XNOR2xp5_ASAP7_75t_R n_5518 (.A(_01000_),
    .B(n_3112_o_0),
    .Y(n_5518_o_0));
 NOR2xp33_ASAP7_75t_R n_5519 (.A(n_5518_o_0),
    .B(n_5517_o_0),
    .Y(n_5519_o_0));
 NOR2xp33_ASAP7_75t_R n_5520 (.A(_00657_),
    .B(net39),
    .Y(n_5520_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5521 (.A1(n_5517_o_0),
    .A2(n_5518_o_0),
    .B(n_5519_o_0),
    .C(net39),
    .D(n_5520_o_0),
    .Y(n_5521_o_0));
 NAND2xp33_ASAP7_75t_R n_5522 (.A(_00880_),
    .B(n_5521_o_0),
    .Y(n_5522_o_0));
 OAI21xp5_ASAP7_75t_R n_5523 (.A1(_00880_),
    .A2(n_5521_o_0),
    .B(n_5522_o_0),
    .Y(n_5523_o_0));
 INVx1_ASAP7_75t_R n_5524 (.A(n_5523_o_0),
    .Y(n_5524_o_0));
 AOI211xp5_ASAP7_75t_R n_5525 (.A1(n_5497_o_0),
    .A2(net39),
    .B(n_5512_o_0),
    .C(n_5498_o_0),
    .Y(n_5525_o_0));
 AOI21x1_ASAP7_75t_R n_5526 (.A1(n_5512_o_0),
    .A2(n_5499_o_0),
    .B(n_5525_o_0),
    .Y(n_5526_o_0));
 INVx1_ASAP7_75t_R n_5527 (.A(n_5490_o_0),
    .Y(n_5527_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5528 (.A1(n_5446_o_0),
    .A2(n_5447_o_0),
    .B(n_5455_o_0),
    .C(net),
    .Y(n_5528_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5529 (.A1(_00529_),
    .A2(net39),
    .B(n_5528_o_0),
    .C(_00877_),
    .Y(n_5529_o_0));
 AOI211xp5_ASAP7_75t_R n_5530 (.A1(_00877_),
    .A2(n_5457_o_0),
    .B(n_5484_o_0),
    .C(n_5529_o_0),
    .Y(n_5530_o_0));
 OAI21xp33_ASAP7_75t_R n_5531 (.A1(n_5530_o_0),
    .A2(n_5489_o_0),
    .B(n_5501_o_0),
    .Y(n_5531_o_0));
 OAI21xp33_ASAP7_75t_R n_5532 (.A1(n_5526_o_0),
    .A2(n_5527_o_0),
    .B(n_5531_o_0),
    .Y(n_5532_o_0));
 NAND2xp33_ASAP7_75t_R n_5533 (.A(_00881_),
    .B(n_5509_o_0),
    .Y(n_5533_o_0));
 OAI21xp33_ASAP7_75t_R n_5534 (.A1(_00881_),
    .A2(n_5509_o_0),
    .B(n_5533_o_0),
    .Y(n_5534_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5535 (.A1(n_5459_o_0),
    .A2(n_5490_o_0),
    .B(n_5532_o_0),
    .C(n_5534_o_0),
    .Y(n_5535_o_0));
 AOI211xp5_ASAP7_75t_R n_5536 (.A1(n_5511_o_0),
    .A2(n_5515_o_0),
    .B(n_5524_o_0),
    .C(n_5535_o_0),
    .Y(n_5536_o_0));
 OAI21xp33_ASAP7_75t_R n_5537 (.A1(n_5483_o_0),
    .A2(n_5459_o_0),
    .B(n_5489_o_0),
    .Y(n_5537_o_0));
 OAI211xp5_ASAP7_75t_R n_5538 (.A1(_00877_),
    .A2(n_5457_o_0),
    .B(n_5484_o_0),
    .C(n_5458_o_0),
    .Y(n_5538_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5539 (.A1(_00877_),
    .A2(n_5457_o_0),
    .B(n_5529_o_0),
    .C(n_5483_o_0),
    .Y(n_5539_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5540 (.A1(n_5538_o_0),
    .A2(n_5539_o_0),
    .B(n_5489_o_0),
    .C(n_5526_o_0),
    .Y(n_5540_o_0));
 INVx1_ASAP7_75t_R n_5541 (.A(n_5540_o_0),
    .Y(n_5541_o_0));
 AOI21xp33_ASAP7_75t_R n_5542 (.A1(n_5537_o_0),
    .A2(n_5541_o_0),
    .B(n_5534_o_0),
    .Y(n_5542_o_0));
 NOR2xp33_ASAP7_75t_R n_5543 (.A(n_5484_o_0),
    .B(n_5459_o_0),
    .Y(n_5543_o_0));
 INVx1_ASAP7_75t_R n_5544 (.A(n_5543_o_0),
    .Y(n_5544_o_0));
 INVx1_ASAP7_75t_R n_5545 (.A(n_5469_o_0),
    .Y(n_5545_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5546 (.A1(_00878_),
    .A2(n_5466_o_0),
    .B(n_5545_o_0),
    .C(n_5484_o_0),
    .Y(n_5546_o_0));
 INVx1_ASAP7_75t_R n_5547 (.A(n_5546_o_0),
    .Y(n_5547_o_0));
 NAND3xp33_ASAP7_75t_R n_5548 (.A(n_5544_o_0),
    .B(n_5547_o_0),
    .C(n_5514_o_0),
    .Y(n_5548_o_0));
 AOI21xp5_ASAP7_75t_R n_5549 (.A1(_00877_),
    .A2(n_5457_o_0),
    .B(n_5529_o_0),
    .Y(n_5549_o_0));
 NOR2xp33_ASAP7_75t_R n_5550 (.A(n_5489_o_0),
    .B(n_5549_o_0),
    .Y(n_5550_o_0));
 INVx1_ASAP7_75t_R n_5551 (.A(n_5550_o_0),
    .Y(n_5551_o_0));
 OAI21xp33_ASAP7_75t_R n_5552 (.A1(n_5459_o_0),
    .A2(n_5490_o_0),
    .B(n_5514_o_0),
    .Y(n_5552_o_0));
 INVx1_ASAP7_75t_R n_5553 (.A(n_5552_o_0),
    .Y(n_5553_o_0));
 AOI21xp33_ASAP7_75t_R n_5554 (.A1(n_5484_o_0),
    .A2(n_5549_o_0),
    .B(n_5489_o_0),
    .Y(n_5554_o_0));
 INVx1_ASAP7_75t_R n_5555 (.A(n_5510_o_0),
    .Y(n_5555_o_0));
 OAI21xp33_ASAP7_75t_R n_5556 (.A1(n_5554_o_0),
    .A2(n_5502_o_0),
    .B(n_5555_o_0),
    .Y(n_5556_o_0));
 XNOR2xp5_ASAP7_75t_R n_5557 (.A(_00880_),
    .B(n_5521_o_0),
    .Y(n_5557_o_0));
 INVx1_ASAP7_75t_R n_5558 (.A(n_5557_o_0),
    .Y(n_5558_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5559 (.A1(n_5551_o_0),
    .A2(n_5553_o_0),
    .B(n_5556_o_0),
    .C(n_5558_o_0),
    .Y(n_5559_o_0));
 AOI21xp33_ASAP7_75t_R n_5560 (.A1(n_5542_o_0),
    .A2(n_5548_o_0),
    .B(n_5559_o_0),
    .Y(n_5560_o_0));
 XNOR2xp5_ASAP7_75t_R n_5561 (.A(_01081_),
    .B(_01082_),
    .Y(n_5561_o_0));
 XNOR2xp5_ASAP7_75t_R n_5562 (.A(_01121_),
    .B(n_5561_o_0),
    .Y(n_5562_o_0));
 XOR2xp5_ASAP7_75t_R n_5563 (.A(_01002_),
    .B(_01041_),
    .Y(n_5563_o_0));
 NOR2xp33_ASAP7_75t_R n_5564 (.A(n_5563_o_0),
    .B(n_5562_o_0),
    .Y(n_5564_o_0));
 NOR2xp33_ASAP7_75t_R n_5565 (.A(_00655_),
    .B(net),
    .Y(n_5565_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5566 (.A1(n_5562_o_0),
    .A2(n_5563_o_0),
    .B(n_5564_o_0),
    .C(net),
    .D(n_5565_o_0),
    .Y(n_5566_o_0));
 XNOR2xp5_ASAP7_75t_R n_5567 (.A(_00882_),
    .B(n_5566_o_0),
    .Y(n_5567_o_0));
 INVx1_ASAP7_75t_R n_5568 (.A(n_5567_o_0),
    .Y(n_5568_o_0));
 OAI21xp33_ASAP7_75t_R n_5569 (.A1(n_5536_o_0),
    .A2(n_5560_o_0),
    .B(n_5568_o_0),
    .Y(n_5569_o_0));
 AOI211xp5_ASAP7_75t_R n_5570 (.A1(n_5497_o_0),
    .A2(net39),
    .B(_00879_),
    .C(n_5498_o_0),
    .Y(n_5570_o_0));
 AOI21x1_ASAP7_75t_R n_5571 (.A1(_00879_),
    .A2(n_5499_o_0),
    .B(n_5570_o_0),
    .Y(n_5571_o_0));
 INVx1_ASAP7_75t_R n_5572 (.A(n_5489_o_0),
    .Y(n_5572_o_0));
 AND2x2_ASAP7_75t_R n_5573 (.A(_00877_),
    .B(n_5457_o_0),
    .Y(n_5573_o_0));
 OAI21xp33_ASAP7_75t_R n_5574 (.A1(n_5529_o_0),
    .A2(n_5573_o_0),
    .B(n_5483_o_0),
    .Y(n_5574_o_0));
 NOR2xp33_ASAP7_75t_R n_5575 (.A(n_5572_o_0),
    .B(n_5574_o_0),
    .Y(n_5575_o_0));
 OAI21xp33_ASAP7_75t_R n_5576 (.A1(n_5529_o_0),
    .A2(n_5573_o_0),
    .B(n_5484_o_0),
    .Y(n_5576_o_0));
 NOR2xp33_ASAP7_75t_R n_5577 (.A(n_5489_o_0),
    .B(n_5576_o_0),
    .Y(n_5577_o_0));
 NAND2xp33_ASAP7_75t_R n_5578 (.A(n_5484_o_0),
    .B(n_5489_o_0),
    .Y(n_5578_o_0));
 INVx1_ASAP7_75t_R n_5579 (.A(n_5578_o_0),
    .Y(n_5579_o_0));
 AOI211xp5_ASAP7_75t_R n_5580 (.A1(_00877_),
    .A2(n_5457_o_0),
    .B(n_5529_o_0),
    .C(n_5483_o_0),
    .Y(n_5580_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5581 (.A1(_00876_),
    .A2(n_5478_o_0),
    .B(n_5482_o_0),
    .C(n_5459_o_0),
    .D(n_5580_o_0),
    .Y(n_5581_o_0));
 OAI21xp33_ASAP7_75t_R n_5582 (.A1(n_5489_o_0),
    .A2(n_5581_o_0),
    .B(n_5571_o_0),
    .Y(n_5582_o_0));
 AO21x1_ASAP7_75t_R n_5583 (.A1(n_5549_o_0),
    .A2(n_5579_o_0),
    .B(n_5582_o_0),
    .Y(n_5583_o_0));
 OAI31xp33_ASAP7_75t_R n_5584 (.A1(n_5571_o_0),
    .A2(n_5575_o_0),
    .A3(n_5577_o_0),
    .B(n_5583_o_0),
    .Y(n_5584_o_0));
 NOR2xp33_ASAP7_75t_R n_5585 (.A(n_5484_o_0),
    .B(n_5549_o_0),
    .Y(n_5585_o_0));
 OAI21xp33_ASAP7_75t_R n_5586 (.A1(n_5489_o_0),
    .A2(n_5483_o_0),
    .B(n_5514_o_0),
    .Y(n_5586_o_0));
 NOR2xp33_ASAP7_75t_R n_5587 (.A(n_5585_o_0),
    .B(n_5586_o_0),
    .Y(n_5587_o_0));
 AOI31xp33_ASAP7_75t_R n_5588 (.A1(n_5501_o_0),
    .A2(n_5578_o_0),
    .A3(n_5544_o_0),
    .B(n_5587_o_0),
    .Y(n_5588_o_0));
 INVx1_ASAP7_75t_R n_5589 (.A(n_5534_o_0),
    .Y(n_5589_o_0));
 OAI21xp33_ASAP7_75t_R n_5590 (.A1(n_5557_o_0),
    .A2(n_5588_o_0),
    .B(n_5589_o_0),
    .Y(n_5590_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5591 (.A1(n_5512_o_0),
    .A2(n_5499_o_0),
    .B(n_5513_o_0),
    .C(n_5489_o_0),
    .Y(n_5591_o_0));
 NAND3xp33_ASAP7_75t_R n_5592 (.A(n_5514_o_0),
    .B(n_5576_o_0),
    .C(net54),
    .Y(n_5592_o_0));
 OAI21xp33_ASAP7_75t_R n_5593 (.A1(n_5540_o_0),
    .A2(n_5575_o_0),
    .B(n_5592_o_0),
    .Y(n_5593_o_0));
 AOI21xp33_ASAP7_75t_R n_5594 (.A1(n_5591_o_0),
    .A2(n_5574_o_0),
    .B(n_5593_o_0),
    .Y(n_5594_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5595 (.A1(n_5572_o_0),
    .A2(n_5581_o_0),
    .B(n_5526_o_0),
    .C(n_5557_o_0),
    .Y(n_5595_o_0));
 NAND2xp33_ASAP7_75t_R n_5596 (.A(n_5489_o_0),
    .B(n_5549_o_0),
    .Y(n_5596_o_0));
 AOI21xp33_ASAP7_75t_R n_5597 (.A1(n_5572_o_0),
    .A2(n_5581_o_0),
    .B(n_5526_o_0),
    .Y(n_5597_o_0));
 NAND2xp33_ASAP7_75t_R n_5598 (.A(n_5596_o_0),
    .B(n_5597_o_0),
    .Y(n_5598_o_0));
 AOI21xp33_ASAP7_75t_R n_5599 (.A1(n_5595_o_0),
    .A2(n_5598_o_0),
    .B(n_5510_o_0),
    .Y(n_5599_o_0));
 NAND2xp33_ASAP7_75t_R n_5600 (.A(_00882_),
    .B(n_5566_o_0),
    .Y(n_5600_o_0));
 OAI21xp33_ASAP7_75t_R n_5601 (.A1(_00882_),
    .A2(n_5566_o_0),
    .B(n_5600_o_0),
    .Y(n_5601_o_0));
 INVx1_ASAP7_75t_R n_5602 (.A(n_5601_o_0),
    .Y(n_5602_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5603 (.A1(n_5524_o_0),
    .A2(n_5594_o_0),
    .B(n_5599_o_0),
    .C(n_5602_o_0),
    .Y(n_5603_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5604 (.A1(n_5523_o_0),
    .A2(n_5584_o_0),
    .B(n_5590_o_0),
    .C(n_5603_o_0),
    .Y(n_5604_o_0));
 OAI31xp33_ASAP7_75t_R n_5605 (.A1(n_5572_o_0),
    .A2(n_5501_o_0),
    .A3(n_5574_o_0),
    .B(n_5523_o_0),
    .Y(n_5605_o_0));
 NAND2xp33_ASAP7_75t_R n_5606 (.A(n_5572_o_0),
    .B(n_5574_o_0),
    .Y(n_5606_o_0));
 AOI21xp33_ASAP7_75t_R n_5607 (.A1(n_5578_o_0),
    .A2(n_5606_o_0),
    .B(n_5514_o_0),
    .Y(n_5607_o_0));
 NOR2xp33_ASAP7_75t_R n_5608 (.A(n_5605_o_0),
    .B(n_5607_o_0),
    .Y(n_5608_o_0));
 INVx1_ASAP7_75t_R n_5609 (.A(n_5530_o_0),
    .Y(n_5609_o_0));
 NOR3xp33_ASAP7_75t_R n_5610 (.A(n_5459_o_0),
    .B(n_5489_o_0),
    .C(n_5484_o_0),
    .Y(n_5610_o_0));
 AOI211xp5_ASAP7_75t_R n_5611 (.A1(n_5609_o_0),
    .A2(n_5489_o_0),
    .B(n_5526_o_0),
    .C(n_5610_o_0),
    .Y(n_5611_o_0));
 INVx1_ASAP7_75t_R n_5612 (.A(n_5611_o_0),
    .Y(n_5612_o_0));
 NOR2xp33_ASAP7_75t_R n_5613 (.A(n_5489_o_0),
    .B(n_5459_o_0),
    .Y(n_5613_o_0));
 AOI31xp33_ASAP7_75t_R n_5614 (.A1(net54),
    .A2(net78),
    .A3(n_5571_o_0),
    .B(n_5557_o_0),
    .Y(n_5614_o_0));
 INVx1_ASAP7_75t_R n_5615 (.A(n_5614_o_0),
    .Y(n_5615_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5616 (.A1(n_5526_o_0),
    .A2(n_5613_o_0),
    .B(n_5615_o_0),
    .C(n_5534_o_0),
    .Y(n_5616_o_0));
 NAND2xp33_ASAP7_75t_R n_5617 (.A(n_5489_o_0),
    .B(n_5576_o_0),
    .Y(n_5617_o_0));
 NAND2xp33_ASAP7_75t_R n_5618 (.A(n_5501_o_0),
    .B(n_5617_o_0),
    .Y(n_5618_o_0));
 INVx1_ASAP7_75t_R n_5619 (.A(n_5574_o_0),
    .Y(n_5619_o_0));
 NAND2xp33_ASAP7_75t_R n_5620 (.A(n_5591_o_0),
    .B(n_5619_o_0),
    .Y(n_5620_o_0));
 OAI21xp33_ASAP7_75t_R n_5621 (.A1(n_5610_o_0),
    .A2(n_5618_o_0),
    .B(n_5620_o_0),
    .Y(n_5621_o_0));
 NOR2xp33_ASAP7_75t_R n_5622 (.A(n_5484_o_0),
    .B(n_5489_o_0),
    .Y(n_5622_o_0));
 OAI21xp33_ASAP7_75t_R n_5623 (.A1(n_5572_o_0),
    .A2(n_5576_o_0),
    .B(n_5514_o_0),
    .Y(n_5623_o_0));
 AOI31xp33_ASAP7_75t_R n_5624 (.A1(n_5572_o_0),
    .A2(n_5619_o_0),
    .A3(n_5526_o_0),
    .B(n_5557_o_0),
    .Y(n_5624_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5625 (.A1(n_5549_o_0),
    .A2(n_5622_o_0),
    .B(n_5623_o_0),
    .C(n_5624_o_0),
    .D(n_5534_o_0),
    .Y(n_5625_o_0));
 OAI21xp33_ASAP7_75t_R n_5626 (.A1(n_5524_o_0),
    .A2(n_5621_o_0),
    .B(n_5625_o_0),
    .Y(n_5626_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5627 (.A1(n_5608_o_0),
    .A2(n_5612_o_0),
    .B(n_5616_o_0),
    .C(n_5626_o_0),
    .Y(n_5627_o_0));
 NOR2xp33_ASAP7_75t_R n_5628 (.A(n_5489_o_0),
    .B(n_5459_o_0),
    .Y(n_5628_o_0));
 AOI211xp5_ASAP7_75t_R n_5629 (.A1(n_5581_o_0),
    .A2(n_5489_o_0),
    .B(n_5526_o_0),
    .C(n_5628_o_0),
    .Y(n_5629_o_0));
 NOR2xp33_ASAP7_75t_R n_5630 (.A(n_5572_o_0),
    .B(n_5576_o_0),
    .Y(n_5630_o_0));
 NOR3xp33_ASAP7_75t_R n_5631 (.A(n_5630_o_0),
    .B(n_5546_o_0),
    .C(n_5571_o_0),
    .Y(n_5631_o_0));
 OAI311xp33_ASAP7_75t_R n_5632 (.A1(n_5574_o_0),
    .A2(n_5526_o_0),
    .A3(net54),
    .B1(n_5524_o_0),
    .C1(n_5531_o_0),
    .Y(n_5632_o_0));
 NOR3xp33_ASAP7_75t_R n_5633 (.A(n_5619_o_0),
    .B(net7),
    .C(n_5526_o_0),
    .Y(n_5633_o_0));
 OAI32xp33_ASAP7_75t_R n_5634 (.A1(n_5629_o_0),
    .A2(n_5631_o_0),
    .A3(n_5558_o_0),
    .B1(n_5632_o_0),
    .B2(n_5633_o_0),
    .Y(n_5634_o_0));
 OAI21xp33_ASAP7_75t_R n_5635 (.A1(n_5555_o_0),
    .A2(n_5634_o_0),
    .B(n_5602_o_0),
    .Y(n_5635_o_0));
 NOR2xp33_ASAP7_75t_R n_5636 (.A(n_5572_o_0),
    .B(n_5526_o_0),
    .Y(n_5636_o_0));
 NAND2xp33_ASAP7_75t_R n_5637 (.A(n_5530_o_0),
    .B(n_5636_o_0),
    .Y(n_5637_o_0));
 OAI31xp33_ASAP7_75t_R n_5638 (.A1(n_5501_o_0),
    .A2(net54),
    .A3(n_5576_o_0),
    .B(n_5558_o_0),
    .Y(n_5638_o_0));
 OAI21xp33_ASAP7_75t_R n_5639 (.A1(n_5486_o_0),
    .A2(n_5502_o_0),
    .B(n_5557_o_0),
    .Y(n_5639_o_0));
 OAI21xp33_ASAP7_75t_R n_5640 (.A1(n_5541_o_0),
    .A2(n_5638_o_0),
    .B(n_5639_o_0),
    .Y(n_5640_o_0));
 AOI21xp33_ASAP7_75t_R n_5641 (.A1(n_5637_o_0),
    .A2(n_5640_o_0),
    .B(n_5589_o_0),
    .Y(n_5641_o_0));
 OAI22xp33_ASAP7_75t_R n_5642 (.A1(n_5627_o_0),
    .A2(n_5568_o_0),
    .B1(n_5635_o_0),
    .B2(n_5641_o_0),
    .Y(n_5642_o_0));
 NOR2xp33_ASAP7_75t_R n_5643 (.A(_00883_),
    .B(n_5442_o_0),
    .Y(n_5643_o_0));
 AND2x2_ASAP7_75t_R n_5644 (.A(_00883_),
    .B(n_5442_o_0),
    .Y(n_5644_o_0));
 NOR2xp33_ASAP7_75t_R n_5645 (.A(n_5643_o_0),
    .B(n_5644_o_0),
    .Y(n_5645_o_0));
 AOI32xp33_ASAP7_75t_R n_5646 (.A1(n_5443_o_0),
    .A2(n_5569_o_0),
    .A3(n_5604_o_0),
    .B1(n_5642_o_0),
    .B2(n_5645_o_0),
    .Y(n_5646_o_0));
 INVx1_ASAP7_75t_R n_5647 (.A(n_5443_o_0),
    .Y(n_5647_o_0));
 OAI221xp5_ASAP7_75t_R n_5648 (.A1(n_5459_o_0),
    .A2(n_5485_o_0),
    .B1(n_5572_o_0),
    .B2(n_5576_o_0),
    .C(n_5514_o_0),
    .Y(n_5648_o_0));
 OAI211xp5_ASAP7_75t_R n_5649 (.A1(net10),
    .A2(n_5549_o_0),
    .B(n_5534_o_0),
    .C(n_5501_o_0),
    .Y(n_5649_o_0));
 OA21x2_ASAP7_75t_R n_5650 (.A1(n_5575_o_0),
    .A2(n_5586_o_0),
    .B(n_5589_o_0),
    .Y(n_5650_o_0));
 OAI211xp5_ASAP7_75t_R n_5651 (.A1(n_5489_o_0),
    .A2(n_5483_o_0),
    .B(n_5501_o_0),
    .C(n_5549_o_0),
    .Y(n_5651_o_0));
 OAI31xp33_ASAP7_75t_R n_5652 (.A1(n_5526_o_0),
    .A2(n_5527_o_0),
    .A3(n_5486_o_0),
    .B(n_5540_o_0),
    .Y(n_5652_o_0));
 OAI21xp33_ASAP7_75t_R n_5653 (.A1(n_5510_o_0),
    .A2(n_5652_o_0),
    .B(n_5568_o_0),
    .Y(n_5653_o_0));
 AO21x1_ASAP7_75t_R n_5654 (.A1(n_5650_o_0),
    .A2(n_5651_o_0),
    .B(n_5653_o_0),
    .Y(n_5654_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5655 (.A1(n_5648_o_0),
    .A2(n_5649_o_0),
    .B(n_5602_o_0),
    .C(n_5654_o_0),
    .Y(n_5655_o_0));
 NOR2xp33_ASAP7_75t_R n_5656 (.A(n_5647_o_0),
    .B(n_5655_o_0),
    .Y(n_5656_o_0));
 INVx1_ASAP7_75t_R n_5657 (.A(n_5645_o_0),
    .Y(n_5657_o_0));
 NOR2xp33_ASAP7_75t_R n_5658 (.A(n_5459_o_0),
    .B(n_5578_o_0),
    .Y(n_5658_o_0));
 OAI21xp33_ASAP7_75t_R n_5659 (.A1(n_5483_o_0),
    .A2(n_5459_o_0),
    .B(n_5539_o_0),
    .Y(n_5659_o_0));
 OAI21xp33_ASAP7_75t_R n_5660 (.A1(n_5489_o_0),
    .A2(n_5659_o_0),
    .B(n_5501_o_0),
    .Y(n_5660_o_0));
 OAI21xp33_ASAP7_75t_R n_5661 (.A1(n_5658_o_0),
    .A2(n_5660_o_0),
    .B(n_5589_o_0),
    .Y(n_5661_o_0));
 AOI31xp33_ASAP7_75t_R n_5662 (.A1(n_5514_o_0),
    .A2(n_5530_o_0),
    .A3(net10),
    .B(n_5661_o_0),
    .Y(n_5662_o_0));
 AOI31xp33_ASAP7_75t_R n_5663 (.A1(n_5539_o_0),
    .A2(n_5538_o_0),
    .A3(n_5489_o_0),
    .B(n_5546_o_0),
    .Y(n_5663_o_0));
 AOI21xp33_ASAP7_75t_R n_5664 (.A1(n_5484_o_0),
    .A2(n_5459_o_0),
    .B(n_5502_o_0),
    .Y(n_5664_o_0));
 AOI211xp5_ASAP7_75t_R n_5665 (.A1(n_5514_o_0),
    .A2(n_5663_o_0),
    .B(n_5664_o_0),
    .C(n_5510_o_0),
    .Y(n_5665_o_0));
 AOI21xp33_ASAP7_75t_R n_5666 (.A1(n_5539_o_0),
    .A2(n_5538_o_0),
    .B(n_5572_o_0),
    .Y(n_5666_o_0));
 NOR3xp33_ASAP7_75t_R n_5667 (.A(n_5666_o_0),
    .B(n_5554_o_0),
    .C(n_5571_o_0),
    .Y(n_5667_o_0));
 AOI21xp33_ASAP7_75t_R n_5668 (.A1(n_5483_o_0),
    .A2(n_5549_o_0),
    .B(n_5571_o_0),
    .Y(n_5668_o_0));
 AO21x1_ASAP7_75t_R n_5669 (.A1(n_5668_o_0),
    .A2(net54),
    .B(n_5534_o_0),
    .Y(n_5669_o_0));
 NOR3xp33_ASAP7_75t_R n_5670 (.A(n_5585_o_0),
    .B(n_5628_o_0),
    .C(n_5526_o_0),
    .Y(n_5670_o_0));
 OAI321xp33_ASAP7_75t_R n_5671 (.A1(n_5510_o_0),
    .A2(n_5611_o_0),
    .A3(n_5667_o_0),
    .B1(n_5669_o_0),
    .B2(n_5670_o_0),
    .C(n_5601_o_0),
    .Y(n_5671_o_0));
 OAI31xp33_ASAP7_75t_R n_5672 (.A1(n_5567_o_0),
    .A2(n_5662_o_0),
    .A3(n_5665_o_0),
    .B(n_5671_o_0),
    .Y(n_5672_o_0));
 OAI21xp33_ASAP7_75t_R n_5673 (.A1(n_5657_o_0),
    .A2(n_5672_o_0),
    .B(n_5523_o_0),
    .Y(n_5673_o_0));
 INVx1_ASAP7_75t_R n_5674 (.A(n_5554_o_0),
    .Y(n_5674_o_0));
 AOI21xp33_ASAP7_75t_R n_5675 (.A1(n_5489_o_0),
    .A2(n_5574_o_0),
    .B(n_5526_o_0),
    .Y(n_5675_o_0));
 AOI21xp33_ASAP7_75t_R n_5676 (.A1(n_5674_o_0),
    .A2(n_5675_o_0),
    .B(n_5510_o_0),
    .Y(n_5676_o_0));
 OA21x2_ASAP7_75t_R n_5677 (.A1(n_5660_o_0),
    .A2(n_5658_o_0),
    .B(n_5676_o_0),
    .Y(n_5677_o_0));
 NAND3xp33_ASAP7_75t_R n_5678 (.A(net78),
    .B(n_5526_o_0),
    .C(net54),
    .Y(n_5678_o_0));
 NAND3xp33_ASAP7_75t_R n_5679 (.A(n_5501_o_0),
    .B(n_5574_o_0),
    .C(net7),
    .Y(n_5679_o_0));
 NAND3xp33_ASAP7_75t_R n_5680 (.A(n_5620_o_0),
    .B(n_5678_o_0),
    .C(n_5679_o_0),
    .Y(n_5680_o_0));
 AOI211xp5_ASAP7_75t_R n_5681 (.A1(n_5514_o_0),
    .A2(n_5579_o_0),
    .B(n_5680_o_0),
    .C(n_5534_o_0),
    .Y(n_5681_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5682 (.A1(n_5549_o_0),
    .A2(net54),
    .B(n_5484_o_0),
    .C(n_5514_o_0),
    .Y(n_5682_o_0));
 INVx1_ASAP7_75t_R n_5683 (.A(n_5682_o_0),
    .Y(n_5683_o_0));
 AOI211xp5_ASAP7_75t_R n_5684 (.A1(n_5484_o_0),
    .A2(n_5549_o_0),
    .B(n_5571_o_0),
    .C(net54),
    .Y(n_5684_o_0));
 INVx1_ASAP7_75t_R n_5685 (.A(n_5596_o_0),
    .Y(n_5685_o_0));
 OA21x2_ASAP7_75t_R n_5686 (.A1(n_5586_o_0),
    .A2(n_5685_o_0),
    .B(n_5555_o_0),
    .Y(n_5686_o_0));
 AOI21xp33_ASAP7_75t_R n_5687 (.A1(n_5651_o_0),
    .A2(n_5686_o_0),
    .B(n_5602_o_0),
    .Y(n_5687_o_0));
 OAI31xp33_ASAP7_75t_R n_5688 (.A1(n_5683_o_0),
    .A2(n_5684_o_0),
    .A3(n_5669_o_0),
    .B(n_5687_o_0),
    .Y(n_5688_o_0));
 OAI31xp33_ASAP7_75t_R n_5689 (.A1(n_5567_o_0),
    .A2(n_5677_o_0),
    .A3(n_5681_o_0),
    .B(n_5688_o_0),
    .Y(n_5689_o_0));
 OAI21xp33_ASAP7_75t_R n_5690 (.A1(n_5489_o_0),
    .A2(n_5530_o_0),
    .B(n_5571_o_0),
    .Y(n_5690_o_0));
 OAI21xp33_ASAP7_75t_R n_5691 (.A1(n_5690_o_0),
    .A2(n_5579_o_0),
    .B(n_5589_o_0),
    .Y(n_5691_o_0));
 NOR2xp33_ASAP7_75t_R n_5692 (.A(n_5527_o_0),
    .B(n_5540_o_0),
    .Y(n_5692_o_0));
 OAI21xp33_ASAP7_75t_R n_5693 (.A1(n_5467_o_0),
    .A2(n_5469_o_0),
    .B(n_5459_o_0),
    .Y(n_5693_o_0));
 NAND2xp33_ASAP7_75t_R n_5694 (.A(n_5501_o_0),
    .B(n_5596_o_0),
    .Y(n_5694_o_0));
 NAND4xp25_ASAP7_75t_R n_5695 (.A(n_5637_o_0),
    .B(n_5693_o_0),
    .C(n_5694_o_0),
    .D(n_5555_o_0),
    .Y(n_5695_o_0));
 OAI211xp5_ASAP7_75t_R n_5696 (.A1(n_5691_o_0),
    .A2(n_5692_o_0),
    .B(n_5695_o_0),
    .C(n_5601_o_0),
    .Y(n_5696_o_0));
 NOR3xp33_ASAP7_75t_R n_5697 (.A(n_5572_o_0),
    .B(n_5459_o_0),
    .C(n_5484_o_0),
    .Y(n_5697_o_0));
 NOR2xp33_ASAP7_75t_R n_5698 (.A(n_5540_o_0),
    .B(n_5697_o_0),
    .Y(n_5698_o_0));
 AOI31xp33_ASAP7_75t_R n_5699 (.A1(n_5514_o_0),
    .A2(n_5578_o_0),
    .A3(n_5606_o_0),
    .B(n_5698_o_0),
    .Y(n_5699_o_0));
 OAI311xp33_ASAP7_75t_R n_5700 (.A1(n_5549_o_0),
    .A2(n_5514_o_0),
    .A3(net54),
    .B1(n_5537_o_0),
    .C1(n_5501_o_0),
    .Y(n_5700_o_0));
 OAI211xp5_ASAP7_75t_R n_5701 (.A1(n_5483_o_0),
    .A2(n_5459_o_0),
    .B(n_5591_o_0),
    .C(n_5571_o_0),
    .Y(n_5701_o_0));
 AOI211xp5_ASAP7_75t_R n_5702 (.A1(n_5700_o_0),
    .A2(n_5701_o_0),
    .B(n_5534_o_0),
    .C(n_5567_o_0),
    .Y(n_5702_o_0));
 AOI31xp33_ASAP7_75t_R n_5703 (.A1(n_5534_o_0),
    .A2(n_5699_o_0),
    .A3(n_5568_o_0),
    .B(n_5702_o_0),
    .Y(n_5703_o_0));
 AOI31xp33_ASAP7_75t_R n_5704 (.A1(n_5696_o_0),
    .A2(n_5703_o_0),
    .A3(n_5645_o_0),
    .B(n_5557_o_0),
    .Y(n_5704_o_0));
 OAI21xp33_ASAP7_75t_R n_5705 (.A1(n_5647_o_0),
    .A2(n_5689_o_0),
    .B(n_5704_o_0),
    .Y(n_5705_o_0));
 OAI21xp33_ASAP7_75t_R n_5706 (.A1(n_5656_o_0),
    .A2(n_5673_o_0),
    .B(n_5705_o_0),
    .Y(n_5706_o_0));
 INVx1_ASAP7_75t_R n_5707 (.A(n_5485_o_0),
    .Y(n_5707_o_0));
 OAI21xp33_ASAP7_75t_R n_5708 (.A1(n_5707_o_0),
    .A2(n_5685_o_0),
    .B(n_5526_o_0),
    .Y(n_5708_o_0));
 INVx1_ASAP7_75t_R n_5709 (.A(n_5629_o_0),
    .Y(n_5709_o_0));
 AOI21xp33_ASAP7_75t_R n_5710 (.A1(n_5708_o_0),
    .A2(n_5709_o_0),
    .B(n_5555_o_0),
    .Y(n_5710_o_0));
 OAI21xp33_ASAP7_75t_R n_5711 (.A1(n_5666_o_0),
    .A2(n_5577_o_0),
    .B(n_5526_o_0),
    .Y(n_5711_o_0));
 OAI211xp5_ASAP7_75t_R n_5712 (.A1(n_5483_o_0),
    .A2(net7),
    .B(n_5514_o_0),
    .C(n_5459_o_0),
    .Y(n_5712_o_0));
 AND3x1_ASAP7_75t_R n_5713 (.A(n_5711_o_0),
    .B(n_5712_o_0),
    .C(n_5555_o_0),
    .Y(n_5713_o_0));
 OAI21xp33_ASAP7_75t_R n_5714 (.A1(n_5572_o_0),
    .A2(n_5581_o_0),
    .B(n_5526_o_0),
    .Y(n_5714_o_0));
 AOI21xp33_ASAP7_75t_R n_5715 (.A1(n_5549_o_0),
    .A2(n_5622_o_0),
    .B(n_5714_o_0),
    .Y(n_5715_o_0));
 AOI21xp33_ASAP7_75t_R n_5716 (.A1(n_5571_o_0),
    .A2(n_5613_o_0),
    .B(n_5715_o_0),
    .Y(n_5716_o_0));
 AOI21xp33_ASAP7_75t_R n_5717 (.A1(n_5459_o_0),
    .A2(net54),
    .B(n_5526_o_0),
    .Y(n_5717_o_0));
 NOR2xp33_ASAP7_75t_R n_5718 (.A(n_5484_o_0),
    .B(n_5549_o_0),
    .Y(n_5718_o_0));
 AOI211xp5_ASAP7_75t_R n_5719 (.A1(n_5549_o_0),
    .A2(n_5572_o_0),
    .B(n_5718_o_0),
    .C(n_5514_o_0),
    .Y(n_5719_o_0));
 OAI21xp33_ASAP7_75t_R n_5720 (.A1(n_5717_o_0),
    .A2(n_5719_o_0),
    .B(n_5555_o_0),
    .Y(n_5720_o_0));
 OAI211xp5_ASAP7_75t_R n_5721 (.A1(n_5716_o_0),
    .A2(n_5534_o_0),
    .B(n_5523_o_0),
    .C(n_5720_o_0),
    .Y(n_5721_o_0));
 OAI31xp33_ASAP7_75t_R n_5722 (.A1(n_5557_o_0),
    .A2(n_5710_o_0),
    .A3(n_5713_o_0),
    .B(n_5721_o_0),
    .Y(n_5722_o_0));
 OAI21xp33_ASAP7_75t_R n_5723 (.A1(n_5571_o_0),
    .A2(n_5613_o_0),
    .B(n_5552_o_0),
    .Y(n_5723_o_0));
 INVx1_ASAP7_75t_R n_5724 (.A(n_5723_o_0),
    .Y(n_5724_o_0));
 OAI21xp33_ASAP7_75t_R n_5725 (.A1(n_5530_o_0),
    .A2(net7),
    .B(n_5541_o_0),
    .Y(n_5725_o_0));
 OAI31xp33_ASAP7_75t_R n_5726 (.A1(net54),
    .A2(n_5526_o_0),
    .A3(n_5619_o_0),
    .B(n_5725_o_0),
    .Y(n_5726_o_0));
 AOI21xp33_ASAP7_75t_R n_5727 (.A1(n_5510_o_0),
    .A2(n_5726_o_0),
    .B(n_5558_o_0),
    .Y(n_5727_o_0));
 OAI21xp33_ASAP7_75t_R n_5728 (.A1(n_5589_o_0),
    .A2(n_5724_o_0),
    .B(n_5727_o_0),
    .Y(n_5728_o_0));
 AOI211xp5_ASAP7_75t_R n_5729 (.A1(n_5483_o_0),
    .A2(n_5549_o_0),
    .B(n_5628_o_0),
    .C(n_5571_o_0),
    .Y(n_5729_o_0));
 AOI31xp33_ASAP7_75t_R n_5730 (.A1(n_5549_o_0),
    .A2(net54),
    .A3(n_5571_o_0),
    .B(n_5729_o_0),
    .Y(n_5730_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5731 (.A1(n_5459_o_0),
    .A2(net54),
    .B(n_5483_o_0),
    .C(n_5501_o_0),
    .Y(n_5731_o_0));
 AO21x1_ASAP7_75t_R n_5732 (.A1(n_5648_o_0),
    .A2(n_5731_o_0),
    .B(n_5555_o_0),
    .Y(n_5732_o_0));
 OAI211xp5_ASAP7_75t_R n_5733 (.A1(n_5730_o_0),
    .A2(n_5510_o_0),
    .B(n_5558_o_0),
    .C(n_5732_o_0),
    .Y(n_5733_o_0));
 AOI31xp33_ASAP7_75t_R n_5734 (.A1(n_5567_o_0),
    .A2(n_5728_o_0),
    .A3(n_5733_o_0),
    .B(n_5443_o_0),
    .Y(n_5734_o_0));
 AOI21xp33_ASAP7_75t_R n_5735 (.A1(n_5549_o_0),
    .A2(n_5526_o_0),
    .B(net54),
    .Y(n_5735_o_0));
 OAI21xp33_ASAP7_75t_R n_5736 (.A1(net10),
    .A2(n_5530_o_0),
    .B(n_5557_o_0),
    .Y(n_5736_o_0));
 NOR2xp33_ASAP7_75t_R n_5737 (.A(n_5483_o_0),
    .B(n_5459_o_0),
    .Y(n_5737_o_0));
 AOI21xp33_ASAP7_75t_R n_5738 (.A1(n_5489_o_0),
    .A2(n_5737_o_0),
    .B(n_5526_o_0),
    .Y(n_5738_o_0));
 OAI32xp33_ASAP7_75t_R n_5739 (.A1(n_5576_o_0),
    .A2(n_5501_o_0),
    .A3(net54),
    .B1(n_5738_o_0),
    .B2(n_5523_o_0),
    .Y(n_5739_o_0));
 OAI31xp33_ASAP7_75t_R n_5740 (.A1(n_5571_o_0),
    .A2(n_5707_o_0),
    .A3(n_5697_o_0),
    .B(n_5739_o_0),
    .Y(n_5740_o_0));
 OAI211xp5_ASAP7_75t_R n_5741 (.A1(n_5735_o_0),
    .A2(n_5736_o_0),
    .B(n_5740_o_0),
    .C(n_5534_o_0),
    .Y(n_5741_o_0));
 AO21x1_ASAP7_75t_R n_5742 (.A1(n_5738_o_0),
    .A2(n_5485_o_0),
    .B(n_5523_o_0),
    .Y(n_5742_o_0));
 NAND2xp33_ASAP7_75t_R n_5743 (.A(n_5489_o_0),
    .B(n_5459_o_0),
    .Y(n_5743_o_0));
 INVx1_ASAP7_75t_R n_5744 (.A(n_5743_o_0),
    .Y(n_5744_o_0));
 NOR3xp33_ASAP7_75t_R n_5745 (.A(n_5577_o_0),
    .B(n_5744_o_0),
    .C(n_5571_o_0),
    .Y(n_5745_o_0));
 OA21x2_ASAP7_75t_R n_5746 (.A1(n_5630_o_0),
    .A2(n_5586_o_0),
    .B(n_5557_o_0),
    .Y(n_5746_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5747 (.A1(n_5660_o_0),
    .A2(n_5666_o_0),
    .B(n_5746_o_0),
    .C(n_5555_o_0),
    .Y(n_5747_o_0));
 OAI21xp33_ASAP7_75t_R n_5748 (.A1(n_5742_o_0),
    .A2(n_5745_o_0),
    .B(n_5747_o_0),
    .Y(n_5748_o_0));
 INVx1_ASAP7_75t_R n_5749 (.A(n_5690_o_0),
    .Y(n_5749_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5750 (.A1(net10),
    .A2(n_5737_o_0),
    .B(n_5749_o_0),
    .C(n_5729_o_0),
    .Y(n_5750_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5751 (.A1(n_5609_o_0),
    .A2(net54),
    .B(n_5610_o_0),
    .C(n_5526_o_0),
    .Y(n_5751_o_0));
 AOI31xp33_ASAP7_75t_R n_5752 (.A1(n_5557_o_0),
    .A2(n_5709_o_0),
    .A3(n_5751_o_0),
    .B(n_5589_o_0),
    .Y(n_5752_o_0));
 AOI21xp33_ASAP7_75t_R n_5753 (.A1(n_5743_o_0),
    .A2(n_5597_o_0),
    .B(n_5523_o_0),
    .Y(n_5753_o_0));
 OAI211xp5_ASAP7_75t_R n_5754 (.A1(n_5574_o_0),
    .A2(n_5572_o_0),
    .B(n_5501_o_0),
    .C(n_5485_o_0),
    .Y(n_5754_o_0));
 OAI221xp5_ASAP7_75t_R n_5755 (.A1(n_5459_o_0),
    .A2(n_5578_o_0),
    .B1(net54),
    .B2(n_5737_o_0),
    .C(n_5501_o_0),
    .Y(n_5755_o_0));
 AOI21xp33_ASAP7_75t_R n_5756 (.A1(n_5552_o_0),
    .A2(n_5755_o_0),
    .B(n_5524_o_0),
    .Y(n_5756_o_0));
 AOI211xp5_ASAP7_75t_R n_5757 (.A1(n_5753_o_0),
    .A2(n_5754_o_0),
    .B(n_5756_o_0),
    .C(n_5555_o_0),
    .Y(n_5757_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5758 (.A1(n_5523_o_0),
    .A2(n_5750_o_0),
    .B(n_5752_o_0),
    .C(n_5757_o_0),
    .Y(n_5758_o_0));
 AOI321xp33_ASAP7_75t_R n_5759 (.A1(n_5602_o_0),
    .A2(n_5741_o_0),
    .A3(n_5748_o_0),
    .B1(n_5758_o_0),
    .B2(n_5567_o_0),
    .C(n_5645_o_0),
    .Y(n_5759_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5760 (.A1(n_5601_o_0),
    .A2(n_5722_o_0),
    .B(n_5734_o_0),
    .C(n_5759_o_0),
    .Y(n_5760_o_0));
 AOI22xp33_ASAP7_75t_R n_5761 (.A1(n_5597_o_0),
    .A2(n_5617_o_0),
    .B1(n_5537_o_0),
    .B2(n_5551_o_0),
    .Y(n_5761_o_0));
 NAND3xp33_ASAP7_75t_R n_5762 (.A(n_5597_o_0),
    .B(n_5617_o_0),
    .C(n_5571_o_0),
    .Y(n_5762_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5763 (.A1(n_5571_o_0),
    .A2(n_5761_o_0),
    .B(n_5762_o_0),
    .C(n_5589_o_0),
    .Y(n_5763_o_0));
 AOI21xp33_ASAP7_75t_R n_5764 (.A1(n_5484_o_0),
    .A2(n_5459_o_0),
    .B(n_5572_o_0),
    .Y(n_5764_o_0));
 OAI21xp33_ASAP7_75t_R n_5765 (.A1(n_5764_o_0),
    .A2(n_5582_o_0),
    .B(n_5589_o_0),
    .Y(n_5765_o_0));
 AOI21xp33_ASAP7_75t_R n_5766 (.A1(n_5578_o_0),
    .A2(n_5668_o_0),
    .B(n_5765_o_0),
    .Y(n_5766_o_0));
 AOI211xp5_ASAP7_75t_R n_5767 (.A1(net10),
    .A2(n_5526_o_0),
    .B(n_5579_o_0),
    .C(n_5585_o_0),
    .Y(n_5767_o_0));
 OA21x2_ASAP7_75t_R n_5768 (.A1(n_5576_o_0),
    .A2(n_5489_o_0),
    .B(n_5490_o_0),
    .Y(n_5768_o_0));
 OAI211xp5_ASAP7_75t_R n_5769 (.A1(n_5549_o_0),
    .A2(net54),
    .B(n_5663_o_0),
    .C(n_5514_o_0),
    .Y(n_5769_o_0));
 OAI31xp33_ASAP7_75t_R n_5770 (.A1(n_5571_o_0),
    .A2(n_5744_o_0),
    .A3(n_5768_o_0),
    .B(n_5769_o_0),
    .Y(n_5770_o_0));
 OAI221xp5_ASAP7_75t_R n_5771 (.A1(n_5510_o_0),
    .A2(n_5767_o_0),
    .B1(n_5534_o_0),
    .B2(n_5770_o_0),
    .C(n_5523_o_0),
    .Y(n_5771_o_0));
 OAI31xp33_ASAP7_75t_R n_5772 (.A1(n_5557_o_0),
    .A2(n_5763_o_0),
    .A3(n_5766_o_0),
    .B(n_5771_o_0),
    .Y(n_5772_o_0));
 NAND2xp33_ASAP7_75t_R n_5773 (.A(net54),
    .B(n_5609_o_0),
    .Y(n_5773_o_0));
 AOI221xp5_ASAP7_75t_R n_5774 (.A1(n_5459_o_0),
    .A2(n_5693_o_0),
    .B1(net7),
    .B2(net78),
    .C(n_5526_o_0),
    .Y(n_5774_o_0));
 AOI31xp33_ASAP7_75t_R n_5775 (.A1(n_5501_o_0),
    .A2(n_5773_o_0),
    .A3(n_5674_o_0),
    .B(n_5774_o_0),
    .Y(n_5775_o_0));
 AOI21xp33_ASAP7_75t_R n_5776 (.A1(n_5483_o_0),
    .A2(n_5459_o_0),
    .B(n_5489_o_0),
    .Y(n_5776_o_0));
 OAI21xp33_ASAP7_75t_R n_5777 (.A1(n_5527_o_0),
    .A2(n_5577_o_0),
    .B(n_5571_o_0),
    .Y(n_5777_o_0));
 OAI211xp5_ASAP7_75t_R n_5778 (.A1(n_5714_o_0),
    .A2(n_5776_o_0),
    .B(n_5777_o_0),
    .C(n_5558_o_0),
    .Y(n_5778_o_0));
 OAI21xp33_ASAP7_75t_R n_5779 (.A1(n_5524_o_0),
    .A2(n_5775_o_0),
    .B(n_5778_o_0),
    .Y(n_5779_o_0));
 OAI21xp33_ASAP7_75t_R n_5780 (.A1(n_5707_o_0),
    .A2(n_5685_o_0),
    .B(n_5571_o_0),
    .Y(n_5780_o_0));
 OAI21xp33_ASAP7_75t_R n_5781 (.A1(n_5543_o_0),
    .A2(n_5586_o_0),
    .B(n_5557_o_0),
    .Y(n_5781_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5782 (.A1(n_5541_o_0),
    .A2(n_5743_o_0),
    .B(n_5781_o_0),
    .C(n_5534_o_0),
    .Y(n_5782_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5783 (.A1(n_5780_o_0),
    .A2(n_5595_o_0),
    .B(n_5782_o_0),
    .C(n_5601_o_0),
    .Y(n_5783_o_0));
 AOI21xp33_ASAP7_75t_R n_5784 (.A1(n_5589_o_0),
    .A2(n_5779_o_0),
    .B(n_5783_o_0),
    .Y(n_5784_o_0));
 AO21x1_ASAP7_75t_R n_5785 (.A1(n_5568_o_0),
    .A2(n_5772_o_0),
    .B(n_5784_o_0),
    .Y(n_5785_o_0));
 OAI21xp33_ASAP7_75t_R n_5786 (.A1(n_5571_o_0),
    .A2(n_5577_o_0),
    .B(n_5746_o_0),
    .Y(n_5786_o_0));
 NOR3xp33_ASAP7_75t_R n_5787 (.A(n_5514_o_0),
    .B(n_5574_o_0),
    .C(net54),
    .Y(n_5787_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5788 (.A1(n_5659_o_0),
    .A2(n_5591_o_0),
    .B(n_5787_o_0),
    .C(n_5524_o_0),
    .Y(n_5788_o_0));
 NAND3xp33_ASAP7_75t_R n_5789 (.A(n_5786_o_0),
    .B(n_5788_o_0),
    .C(n_5510_o_0),
    .Y(n_5789_o_0));
 NOR2xp33_ASAP7_75t_R n_5790 (.A(n_5483_o_0),
    .B(n_5489_o_0),
    .Y(n_5790_o_0));
 INVx1_ASAP7_75t_R n_5791 (.A(n_5790_o_0),
    .Y(n_5791_o_0));
 AOI31xp33_ASAP7_75t_R n_5792 (.A1(n_5501_o_0),
    .A2(n_5791_o_0),
    .A3(n_5537_o_0),
    .B(n_5558_o_0),
    .Y(n_5792_o_0));
 OA21x2_ASAP7_75t_R n_5793 (.A1(n_5527_o_0),
    .A2(n_5582_o_0),
    .B(n_5792_o_0),
    .Y(n_5793_o_0));
 INVx1_ASAP7_75t_R n_5794 (.A(n_5623_o_0),
    .Y(n_5794_o_0));
 OAI31xp33_ASAP7_75t_R n_5795 (.A1(net7),
    .A2(n_5514_o_0),
    .A3(net78),
    .B(n_5624_o_0),
    .Y(n_5795_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5796 (.A1(n_5459_o_0),
    .A2(net54),
    .B(n_5794_o_0),
    .C(n_5795_o_0),
    .Y(n_5796_o_0));
 OAI21xp33_ASAP7_75t_R n_5797 (.A1(n_5793_o_0),
    .A2(n_5796_o_0),
    .B(n_5534_o_0),
    .Y(n_5797_o_0));
 AOI21xp33_ASAP7_75t_R n_5798 (.A1(n_5572_o_0),
    .A2(n_5659_o_0),
    .B(n_5501_o_0),
    .Y(n_5798_o_0));
 NAND3xp33_ASAP7_75t_R n_5799 (.A(n_5572_o_0),
    .B(n_5459_o_0),
    .C(n_5484_o_0),
    .Y(n_5799_o_0));
 AOI21xp33_ASAP7_75t_R n_5800 (.A1(n_5490_o_0),
    .A2(n_5799_o_0),
    .B(n_5514_o_0),
    .Y(n_5800_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5801 (.A1(net10),
    .A2(n_5737_o_0),
    .B(n_5798_o_0),
    .C(n_5800_o_0),
    .Y(n_5801_o_0));
 AOI211xp5_ASAP7_75t_R n_5802 (.A1(n_5549_o_0),
    .A2(net7),
    .B(n_5718_o_0),
    .C(n_5501_o_0),
    .Y(n_5802_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5803 (.A1(n_5802_o_0),
    .A2(n_5607_o_0),
    .B(n_5557_o_0),
    .C(n_5555_o_0),
    .Y(n_5803_o_0));
 OAI31xp33_ASAP7_75t_R n_5804 (.A1(n_5571_o_0),
    .A2(n_5764_o_0),
    .A3(n_5790_o_0),
    .B(n_5648_o_0),
    .Y(n_5804_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5805 (.A1(n_5738_o_0),
    .A2(n_5485_o_0),
    .B(n_5523_o_0),
    .C(n_5534_o_0),
    .Y(n_5805_o_0));
 AOI21xp33_ASAP7_75t_R n_5806 (.A1(n_5557_o_0),
    .A2(n_5804_o_0),
    .B(n_5805_o_0),
    .Y(n_5806_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5807 (.A1(n_5523_o_0),
    .A2(n_5801_o_0),
    .B(n_5803_o_0),
    .C(n_5806_o_0),
    .Y(n_5807_o_0));
 AOI321xp33_ASAP7_75t_R n_5808 (.A1(n_5789_o_0),
    .A2(n_5797_o_0),
    .A3(n_5567_o_0),
    .B1(n_5602_o_0),
    .B2(n_5807_o_0),
    .C(n_5645_o_0),
    .Y(n_5808_o_0));
 AOI21xp33_ASAP7_75t_R n_5809 (.A1(n_5647_o_0),
    .A2(n_5785_o_0),
    .B(n_5808_o_0),
    .Y(n_5809_o_0));
 INVx1_ASAP7_75t_R n_5810 (.A(n_5675_o_0),
    .Y(n_5810_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5811 (.A1(n_5459_o_0),
    .A2(n_5578_o_0),
    .B(n_5501_o_0),
    .C(n_5523_o_0),
    .Y(n_5811_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5812 (.A1(net54),
    .A2(net78),
    .B(n_5690_o_0),
    .C(n_5557_o_0),
    .Y(n_5812_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5813 (.A1(n_5487_o_0),
    .A2(n_5503_o_0),
    .B(n_5812_o_0),
    .C(n_5510_o_0),
    .Y(n_5813_o_0));
 INVx1_ASAP7_75t_R n_5814 (.A(n_5537_o_0),
    .Y(n_5814_o_0));
 AOI21xp33_ASAP7_75t_R n_5815 (.A1(n_5483_o_0),
    .A2(n_5514_o_0),
    .B(net54),
    .Y(n_5815_o_0));
 AOI21xp33_ASAP7_75t_R n_5816 (.A1(n_5571_o_0),
    .A2(n_5814_o_0),
    .B(n_5815_o_0),
    .Y(n_5816_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5817 (.A1(net54),
    .A2(n_5459_o_0),
    .B(n_5776_o_0),
    .C(n_5514_o_0),
    .Y(n_5817_o_0));
 AOI31xp33_ASAP7_75t_R n_5818 (.A1(n_5651_o_0),
    .A2(n_5817_o_0),
    .A3(n_5524_o_0),
    .B(n_5589_o_0),
    .Y(n_5818_o_0));
 OAI21xp33_ASAP7_75t_R n_5819 (.A1(n_5558_o_0),
    .A2(n_5816_o_0),
    .B(n_5818_o_0),
    .Y(n_5819_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5820 (.A1(n_5810_o_0),
    .A2(n_5811_o_0),
    .B(n_5813_o_0),
    .C(n_5819_o_0),
    .Y(n_5820_o_0));
 NOR2xp33_ASAP7_75t_R n_5821 (.A(n_5647_o_0),
    .B(n_5820_o_0),
    .Y(n_5821_o_0));
 NOR2xp33_ASAP7_75t_R n_5822 (.A(n_5586_o_0),
    .B(n_5685_o_0),
    .Y(n_5822_o_0));
 OAI21xp33_ASAP7_75t_R n_5823 (.A1(n_5543_o_0),
    .A2(n_5744_o_0),
    .B(n_5571_o_0),
    .Y(n_5823_o_0));
 OAI311xp33_ASAP7_75t_R n_5824 (.A1(n_5571_o_0),
    .A2(n_5575_o_0),
    .A3(n_5550_o_0),
    .B1(n_5558_o_0),
    .C1(n_5823_o_0),
    .Y(n_5824_o_0));
 OAI31xp33_ASAP7_75t_R n_5825 (.A1(n_5524_o_0),
    .A2(n_5719_o_0),
    .A3(n_5822_o_0),
    .B(n_5824_o_0),
    .Y(n_5825_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5826 (.A1(n_5484_o_0),
    .A2(n_5459_o_0),
    .B(n_5572_o_0),
    .C(n_5526_o_0),
    .Y(n_5826_o_0));
 OAI211xp5_ASAP7_75t_R n_5827 (.A1(n_5574_o_0),
    .A2(net54),
    .B(n_5826_o_0),
    .C(n_5558_o_0),
    .Y(n_5827_o_0));
 NAND2xp33_ASAP7_75t_R n_5828 (.A(n_5596_o_0),
    .B(n_5547_o_0),
    .Y(n_5828_o_0));
 OAI211xp5_ASAP7_75t_R n_5829 (.A1(n_5828_o_0),
    .A2(n_5571_o_0),
    .B(n_5682_o_0),
    .C(n_5557_o_0),
    .Y(n_5829_o_0));
 AOI21xp33_ASAP7_75t_R n_5830 (.A1(n_5827_o_0),
    .A2(n_5829_o_0),
    .B(n_5534_o_0),
    .Y(n_5830_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5831 (.A1(n_5825_o_0),
    .A2(n_5534_o_0),
    .B(n_5830_o_0),
    .C(n_5645_o_0),
    .Y(n_5831_o_0));
 INVx1_ASAP7_75t_R n_5832 (.A(n_5831_o_0),
    .Y(n_5832_o_0));
 OAI21xp33_ASAP7_75t_R n_5833 (.A1(n_5526_o_0),
    .A2(n_5737_o_0),
    .B(n_5557_o_0),
    .Y(n_5833_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5834 (.A1(net10),
    .A2(n_5659_o_0),
    .B(n_5501_o_0),
    .C(n_5833_o_0),
    .Y(n_5834_o_0));
 OAI21xp33_ASAP7_75t_R n_5835 (.A1(n_5550_o_0),
    .A2(n_5618_o_0),
    .B(n_5524_o_0),
    .Y(n_5835_o_0));
 AOI21xp33_ASAP7_75t_R n_5836 (.A1(n_5591_o_0),
    .A2(n_5544_o_0),
    .B(n_5835_o_0),
    .Y(n_5836_o_0));
 OAI21xp33_ASAP7_75t_R n_5837 (.A1(n_5834_o_0),
    .A2(n_5836_o_0),
    .B(n_5589_o_0),
    .Y(n_5837_o_0));
 NAND2xp33_ASAP7_75t_R n_5838 (.A(n_5558_o_0),
    .B(n_5823_o_0),
    .Y(n_5838_o_0));
 AOI22xp33_ASAP7_75t_R n_5839 (.A1(n_5636_o_0),
    .A2(n_5574_o_0),
    .B1(n_5578_o_0),
    .B2(n_5668_o_0),
    .Y(n_5839_o_0));
 OAI31xp33_ASAP7_75t_R n_5840 (.A1(n_5574_o_0),
    .A2(n_5526_o_0),
    .A3(net54),
    .B(n_5839_o_0),
    .Y(n_5840_o_0));
 AOI21xp33_ASAP7_75t_R n_5841 (.A1(n_5523_o_0),
    .A2(n_5840_o_0),
    .B(n_5510_o_0),
    .Y(n_5841_o_0));
 OAI21xp33_ASAP7_75t_R n_5842 (.A1(n_5838_o_0),
    .A2(n_5631_o_0),
    .B(n_5841_o_0),
    .Y(n_5842_o_0));
 INVx1_ASAP7_75t_R n_5843 (.A(n_5610_o_0),
    .Y(n_5843_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5844 (.A1(n_5484_o_0),
    .A2(n_5549_o_0),
    .B(n_5489_o_0),
    .C(n_5571_o_0),
    .Y(n_5844_o_0));
 OAI21xp33_ASAP7_75t_R n_5845 (.A1(n_5666_o_0),
    .A2(n_5844_o_0),
    .B(n_5557_o_0),
    .Y(n_5845_o_0));
 AOI31xp33_ASAP7_75t_R n_5846 (.A1(n_5501_o_0),
    .A2(n_5843_o_0),
    .A3(n_5617_o_0),
    .B(n_5845_o_0),
    .Y(n_5846_o_0));
 OAI31xp33_ASAP7_75t_R n_5847 (.A1(n_5572_o_0),
    .A2(n_5514_o_0),
    .A3(n_5659_o_0),
    .B(n_5799_o_0),
    .Y(n_5847_o_0));
 AOI211xp5_ASAP7_75t_R n_5848 (.A1(n_5530_o_0),
    .A2(n_5636_o_0),
    .B(n_5847_o_0),
    .C(n_5523_o_0),
    .Y(n_5848_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5849 (.A1(net54),
    .A2(n_5483_o_0),
    .B(n_5459_o_0),
    .C(n_5571_o_0),
    .Y(n_5849_o_0));
 OAI211xp5_ASAP7_75t_R n_5850 (.A1(n_5530_o_0),
    .A2(n_5489_o_0),
    .B(n_5537_o_0),
    .C(n_5571_o_0),
    .Y(n_5850_o_0));
 OAI31xp33_ASAP7_75t_R n_5851 (.A1(n_5571_o_0),
    .A2(n_5744_o_0),
    .A3(n_5610_o_0),
    .B(n_5850_o_0),
    .Y(n_5851_o_0));
 OAI321xp33_ASAP7_75t_R n_5852 (.A1(n_5558_o_0),
    .A2(n_5611_o_0),
    .A3(n_5849_o_0),
    .B1(n_5851_o_0),
    .B2(n_5523_o_0),
    .C(n_5534_o_0),
    .Y(n_5852_o_0));
 OAI31xp33_ASAP7_75t_R n_5853 (.A1(n_5555_o_0),
    .A2(n_5846_o_0),
    .A3(n_5848_o_0),
    .B(n_5852_o_0),
    .Y(n_5853_o_0));
 NOR2xp33_ASAP7_75t_R n_5854 (.A(n_5602_o_0),
    .B(n_5645_o_0),
    .Y(n_5854_o_0));
 AO31x2_ASAP7_75t_R n_5855 (.A1(n_5853_o_0),
    .A2(n_5601_o_0),
    .A3(n_5645_o_0),
    .B(n_5854_o_0),
    .Y(n_5855_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5856 (.A1(n_5837_o_0),
    .A2(n_5842_o_0),
    .B(n_5647_o_0),
    .C(n_5855_o_0),
    .Y(n_5856_o_0));
 OAI31xp33_ASAP7_75t_R n_5857 (.A1(n_5567_o_0),
    .A2(n_5821_o_0),
    .A3(n_5832_o_0),
    .B(n_5856_o_0),
    .Y(n_5857_o_0));
 NOR3xp33_ASAP7_75t_R n_5858 (.A(n_5764_o_0),
    .B(n_5610_o_0),
    .C(n_5526_o_0),
    .Y(n_5858_o_0));
 AOI31xp33_ASAP7_75t_R n_5859 (.A1(n_5483_o_0),
    .A2(n_5501_o_0),
    .A3(n_5773_o_0),
    .B(n_5858_o_0),
    .Y(n_5859_o_0));
 OA211x2_ASAP7_75t_R n_5860 (.A1(n_5531_o_0),
    .A2(n_5814_o_0),
    .B(n_5515_o_0),
    .C(n_5557_o_0),
    .Y(n_5860_o_0));
 AOI211xp5_ASAP7_75t_R n_5861 (.A1(n_5859_o_0),
    .A2(n_5524_o_0),
    .B(n_5555_o_0),
    .C(n_5860_o_0),
    .Y(n_5861_o_0));
 NAND4xp25_ASAP7_75t_R n_5862 (.A(n_5690_o_0),
    .B(n_5558_o_0),
    .C(n_5578_o_0),
    .D(n_5743_o_0),
    .Y(n_5862_o_0));
 OAI31xp33_ASAP7_75t_R n_5863 (.A1(n_5524_o_0),
    .A2(n_5798_o_0),
    .A3(n_5800_o_0),
    .B(n_5862_o_0),
    .Y(n_5863_o_0));
 OAI21xp33_ASAP7_75t_R n_5864 (.A1(n_5510_o_0),
    .A2(n_5863_o_0),
    .B(n_5568_o_0),
    .Y(n_5864_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5865 (.A1(net10),
    .A2(n_5619_o_0),
    .B(n_5541_o_0),
    .C(n_5738_o_0),
    .Y(n_5865_o_0));
 OAI211xp5_ASAP7_75t_R n_5866 (.A1(n_5810_o_0),
    .A2(n_5628_o_0),
    .B(n_5678_o_0),
    .C(n_5524_o_0),
    .Y(n_5866_o_0));
 OAI21xp33_ASAP7_75t_R n_5867 (.A1(n_5524_o_0),
    .A2(n_5865_o_0),
    .B(n_5866_o_0),
    .Y(n_5867_o_0));
 OAI21xp33_ASAP7_75t_R n_5868 (.A1(n_5459_o_0),
    .A2(n_5514_o_0),
    .B(n_5823_o_0),
    .Y(n_5868_o_0));
 NOR3xp33_ASAP7_75t_R n_5869 (.A(n_5764_o_0),
    .B(n_5550_o_0),
    .C(n_5546_o_0),
    .Y(n_5869_o_0));
 AOI211xp5_ASAP7_75t_R n_5870 (.A1(n_5484_o_0),
    .A2(n_5549_o_0),
    .B(n_5527_o_0),
    .C(n_5526_o_0),
    .Y(n_5870_o_0));
 AOI211xp5_ASAP7_75t_R n_5871 (.A1(n_5869_o_0),
    .A2(n_5501_o_0),
    .B(n_5870_o_0),
    .C(n_5523_o_0),
    .Y(n_5871_o_0));
 AOI211xp5_ASAP7_75t_R n_5872 (.A1(n_5868_o_0),
    .A2(n_5557_o_0),
    .B(n_5871_o_0),
    .C(n_5555_o_0),
    .Y(n_5872_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5873 (.A1(n_5534_o_0),
    .A2(n_5867_o_0),
    .B(n_5872_o_0),
    .C(n_5567_o_0),
    .Y(n_5873_o_0));
 OAI21xp33_ASAP7_75t_R n_5874 (.A1(n_5861_o_0),
    .A2(n_5864_o_0),
    .B(n_5873_o_0),
    .Y(n_5874_o_0));
 AOI22xp33_ASAP7_75t_R n_5875 (.A1(n_5503_o_0),
    .A2(n_5487_o_0),
    .B1(n_5530_o_0),
    .B2(n_5636_o_0),
    .Y(n_5875_o_0));
 AOI21xp33_ASAP7_75t_R n_5876 (.A1(n_5484_o_0),
    .A2(n_5591_o_0),
    .B(n_5510_o_0),
    .Y(n_5876_o_0));
 OAI21xp33_ASAP7_75t_R n_5877 (.A1(n_5585_o_0),
    .A2(n_5586_o_0),
    .B(n_5589_o_0),
    .Y(n_5877_o_0));
 AOI21xp33_ASAP7_75t_R n_5878 (.A1(n_5484_o_0),
    .A2(n_5501_o_0),
    .B(n_5877_o_0),
    .Y(n_5878_o_0));
 AOI21xp33_ASAP7_75t_R n_5879 (.A1(n_5875_o_0),
    .A2(n_5876_o_0),
    .B(n_5878_o_0),
    .Y(n_5879_o_0));
 AOI211xp5_ASAP7_75t_R n_5880 (.A1(n_5484_o_0),
    .A2(n_5459_o_0),
    .B(n_5571_o_0),
    .C(net7),
    .Y(n_5880_o_0));
 AOI31xp33_ASAP7_75t_R n_5881 (.A1(n_5514_o_0),
    .A2(n_5487_o_0),
    .A3(n_5537_o_0),
    .B(n_5880_o_0),
    .Y(n_5881_o_0));
 OAI221xp5_ASAP7_75t_R n_5882 (.A1(n_5459_o_0),
    .A2(n_5490_o_0),
    .B1(net54),
    .B2(n_5581_o_0),
    .C(n_5526_o_0),
    .Y(n_5882_o_0));
 OAI31xp33_ASAP7_75t_R n_5883 (.A1(n_5526_o_0),
    .A2(n_5764_o_0),
    .A3(n_5550_o_0),
    .B(n_5882_o_0),
    .Y(n_5883_o_0));
 AOI21xp33_ASAP7_75t_R n_5884 (.A1(n_5510_o_0),
    .A2(n_5883_o_0),
    .B(n_5523_o_0),
    .Y(n_5884_o_0));
 OAI21xp33_ASAP7_75t_R n_5885 (.A1(n_5589_o_0),
    .A2(n_5881_o_0),
    .B(n_5884_o_0),
    .Y(n_5885_o_0));
 OAI21xp33_ASAP7_75t_R n_5886 (.A1(n_5558_o_0),
    .A2(n_5879_o_0),
    .B(n_5885_o_0),
    .Y(n_5886_o_0));
 AOI22xp33_ASAP7_75t_R n_5887 (.A1(n_5636_o_0),
    .A2(n_5530_o_0),
    .B1(n_5537_o_0),
    .B2(n_5501_o_0),
    .Y(n_5887_o_0));
 OAI21xp33_ASAP7_75t_R n_5888 (.A1(n_5540_o_0),
    .A2(n_5630_o_0),
    .B(n_5555_o_0),
    .Y(n_5888_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5889 (.A1(n_5537_o_0),
    .A2(n_5597_o_0),
    .B(n_5888_o_0),
    .C(n_5558_o_0),
    .Y(n_5889_o_0));
 NOR2xp33_ASAP7_75t_R n_5890 (.A(_00880_),
    .B(n_5521_o_0),
    .Y(n_5890_o_0));
 INVx1_ASAP7_75t_R n_5891 (.A(n_5522_o_0),
    .Y(n_5891_o_0));
 AOI21xp33_ASAP7_75t_R n_5892 (.A1(n_5576_o_0),
    .A2(n_5501_o_0),
    .B(n_5510_o_0),
    .Y(n_5892_o_0));
 OAI21xp33_ASAP7_75t_R n_5893 (.A1(n_5526_o_0),
    .A2(n_5486_o_0),
    .B(n_5892_o_0),
    .Y(n_5893_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5894 (.A1(n_5483_o_0),
    .A2(net54),
    .B(n_5501_o_0),
    .C(n_5534_o_0),
    .Y(n_5894_o_0));
 OAI21xp33_ASAP7_75t_R n_5895 (.A1(n_5552_o_0),
    .A2(n_5486_o_0),
    .B(n_5894_o_0),
    .Y(n_5895_o_0));
 OAI211xp5_ASAP7_75t_R n_5896 (.A1(n_5890_o_0),
    .A2(n_5891_o_0),
    .B(n_5893_o_0),
    .C(n_5895_o_0),
    .Y(n_5896_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5897 (.A1(n_5589_o_0),
    .A2(n_5887_o_0),
    .B(n_5889_o_0),
    .C(n_5896_o_0),
    .Y(n_5897_o_0));
 OAI22xp33_ASAP7_75t_R n_5898 (.A1(n_5897_o_0),
    .A2(n_5568_o_0),
    .B1(n_5644_o_0),
    .B2(n_5643_o_0),
    .Y(n_5898_o_0));
 AO21x1_ASAP7_75t_R n_5899 (.A1(n_5602_o_0),
    .A2(n_5886_o_0),
    .B(n_5898_o_0),
    .Y(n_5899_o_0));
 OAI21xp33_ASAP7_75t_R n_5900 (.A1(n_5443_o_0),
    .A2(n_5874_o_0),
    .B(n_5899_o_0),
    .Y(n_5900_o_0));
 INVx1_ASAP7_75t_R n_5901 (.A(n_5844_o_0),
    .Y(n_5901_o_0));
 AOI211xp5_ASAP7_75t_R n_5902 (.A1(net10),
    .A2(n_5574_o_0),
    .B(n_5658_o_0),
    .C(n_5571_o_0),
    .Y(n_5902_o_0));
 AOI21xp33_ASAP7_75t_R n_5903 (.A1(n_5901_o_0),
    .A2(n_5617_o_0),
    .B(n_5902_o_0),
    .Y(n_5903_o_0));
 OAI211xp5_ASAP7_75t_R n_5904 (.A1(net7),
    .A2(n_5484_o_0),
    .B(n_5799_o_0),
    .C(n_5501_o_0),
    .Y(n_5904_o_0));
 OAI211xp5_ASAP7_75t_R n_5905 (.A1(n_5501_o_0),
    .A2(n_5485_o_0),
    .B(n_5614_o_0),
    .C(n_5904_o_0),
    .Y(n_5905_o_0));
 OAI21xp33_ASAP7_75t_R n_5906 (.A1(n_5524_o_0),
    .A2(n_5903_o_0),
    .B(n_5905_o_0),
    .Y(n_5906_o_0));
 AOI221xp5_ASAP7_75t_R n_5907 (.A1(n_5459_o_0),
    .A2(n_5571_o_0),
    .B1(n_5743_o_0),
    .B2(n_5668_o_0),
    .C(n_5524_o_0),
    .Y(n_5907_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5908 (.A1(n_5575_o_0),
    .A2(n_5577_o_0),
    .B(n_5526_o_0),
    .C(n_5557_o_0),
    .Y(n_5908_o_0));
 OA21x2_ASAP7_75t_R n_5909 (.A1(n_5501_o_0),
    .A2(n_5606_o_0),
    .B(n_5908_o_0),
    .Y(n_5909_o_0));
 OAI31xp33_ASAP7_75t_R n_5910 (.A1(n_5907_o_0),
    .A2(n_5909_o_0),
    .A3(n_5534_o_0),
    .B(n_5568_o_0),
    .Y(n_5910_o_0));
 AOI21xp33_ASAP7_75t_R n_5911 (.A1(n_5555_o_0),
    .A2(n_5906_o_0),
    .B(n_5910_o_0),
    .Y(n_5911_o_0));
 OAI311xp33_ASAP7_75t_R n_5912 (.A1(net54),
    .A2(n_5526_o_0),
    .A3(net78),
    .B1(n_5558_o_0),
    .C1(n_5723_o_0),
    .Y(n_5912_o_0));
 NOR2xp33_ASAP7_75t_R n_5913 (.A(n_5459_o_0),
    .B(n_5490_o_0),
    .Y(n_5913_o_0));
 OAI21xp33_ASAP7_75t_R n_5914 (.A1(net54),
    .A2(n_5659_o_0),
    .B(n_5675_o_0),
    .Y(n_5914_o_0));
 OAI31xp33_ASAP7_75t_R n_5915 (.A1(n_5571_o_0),
    .A2(n_5913_o_0),
    .A3(n_5550_o_0),
    .B(n_5914_o_0),
    .Y(n_5915_o_0));
 AOI21xp33_ASAP7_75t_R n_5916 (.A1(n_5523_o_0),
    .A2(n_5915_o_0),
    .B(n_5534_o_0),
    .Y(n_5916_o_0));
 OAI211xp5_ASAP7_75t_R n_5917 (.A1(net7),
    .A2(n_5659_o_0),
    .B(n_5791_o_0),
    .C(n_5514_o_0),
    .Y(n_5917_o_0));
 OAI31xp33_ASAP7_75t_R n_5918 (.A1(n_5571_o_0),
    .A2(n_5610_o_0),
    .A3(n_5579_o_0),
    .B(n_5917_o_0),
    .Y(n_5918_o_0));
 AOI22xp33_ASAP7_75t_R n_5919 (.A1(n_5636_o_0),
    .A2(n_5576_o_0),
    .B1(n_5596_o_0),
    .B2(n_5668_o_0),
    .Y(n_5919_o_0));
 OAI21xp33_ASAP7_75t_R n_5920 (.A1(n_5557_o_0),
    .A2(n_5919_o_0),
    .B(n_5555_o_0),
    .Y(n_5920_o_0));
 AOI21xp33_ASAP7_75t_R n_5921 (.A1(n_5523_o_0),
    .A2(n_5918_o_0),
    .B(n_5920_o_0),
    .Y(n_5921_o_0));
 AOI21xp33_ASAP7_75t_R n_5922 (.A1(n_5912_o_0),
    .A2(n_5916_o_0),
    .B(n_5921_o_0),
    .Y(n_5922_o_0));
 OAI21xp33_ASAP7_75t_R n_5923 (.A1(n_5602_o_0),
    .A2(n_5922_o_0),
    .B(n_5645_o_0),
    .Y(n_5923_o_0));
 OAI21xp33_ASAP7_75t_R n_5924 (.A1(n_5707_o_0),
    .A2(n_5543_o_0),
    .B(n_5526_o_0),
    .Y(n_5924_o_0));
 AOI21xp33_ASAP7_75t_R n_5925 (.A1(n_5844_o_0),
    .A2(n_5924_o_0),
    .B(n_5523_o_0),
    .Y(n_5925_o_0));
 OAI21xp33_ASAP7_75t_R n_5926 (.A1(n_5578_o_0),
    .A2(n_5526_o_0),
    .B(n_5925_o_0),
    .Y(n_5926_o_0));
 AOI21xp33_ASAP7_75t_R n_5927 (.A1(n_5484_o_0),
    .A2(n_5501_o_0),
    .B(n_5549_o_0),
    .Y(n_5927_o_0));
 OAI21xp33_ASAP7_75t_R n_5928 (.A1(n_5579_o_0),
    .A2(n_5927_o_0),
    .B(n_5557_o_0),
    .Y(n_5928_o_0));
 AOI21xp33_ASAP7_75t_R n_5929 (.A1(n_5799_o_0),
    .A2(n_5503_o_0),
    .B(n_5597_o_0),
    .Y(n_5929_o_0));
 AOI21xp33_ASAP7_75t_R n_5930 (.A1(n_5501_o_0),
    .A2(n_5596_o_0),
    .B(n_5523_o_0),
    .Y(n_5930_o_0));
 AOI21xp33_ASAP7_75t_R n_5931 (.A1(n_5930_o_0),
    .A2(n_5548_o_0),
    .B(n_5589_o_0),
    .Y(n_5931_o_0));
 OAI21xp33_ASAP7_75t_R n_5932 (.A1(n_5524_o_0),
    .A2(n_5929_o_0),
    .B(n_5931_o_0),
    .Y(n_5932_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5933 (.A1(n_5926_o_0),
    .A2(n_5928_o_0),
    .B(n_5534_o_0),
    .C(n_5932_o_0),
    .Y(n_5933_o_0));
 OAI21xp33_ASAP7_75t_R n_5934 (.A1(n_5814_o_0),
    .A2(n_5660_o_0),
    .B(n_5524_o_0),
    .Y(n_5934_o_0));
 OAI21xp33_ASAP7_75t_R n_5935 (.A1(n_5459_o_0),
    .A2(n_5572_o_0),
    .B(n_5693_o_0),
    .Y(n_5935_o_0));
 OAI31xp33_ASAP7_75t_R n_5936 (.A1(n_5526_o_0),
    .A2(n_5764_o_0),
    .A3(n_5550_o_0),
    .B(n_5557_o_0),
    .Y(n_5936_o_0));
 AO21x1_ASAP7_75t_R n_5937 (.A1(n_5501_o_0),
    .A2(n_5935_o_0),
    .B(n_5936_o_0),
    .Y(n_5937_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5938 (.A1(n_5514_o_0),
    .A2(n_5579_o_0),
    .B(n_5934_o_0),
    .C(n_5937_o_0),
    .Y(n_5938_o_0));
 INVx1_ASAP7_75t_R n_5939 (.A(n_5693_o_0),
    .Y(n_5939_o_0));
 OAI211xp5_ASAP7_75t_R n_5940 (.A1(n_5826_o_0),
    .A2(n_5939_o_0),
    .B(n_5558_o_0),
    .C(n_5623_o_0),
    .Y(n_5940_o_0));
 OAI211xp5_ASAP7_75t_R n_5941 (.A1(n_5524_o_0),
    .A2(n_5751_o_0),
    .B(n_5940_o_0),
    .C(n_5555_o_0),
    .Y(n_5941_o_0));
 OAI211xp5_ASAP7_75t_R n_5942 (.A1(n_5938_o_0),
    .A2(n_5555_o_0),
    .B(n_5567_o_0),
    .C(n_5941_o_0),
    .Y(n_5942_o_0));
 OAI211xp5_ASAP7_75t_R n_5943 (.A1(n_5933_o_0),
    .A2(n_5567_o_0),
    .B(n_5942_o_0),
    .C(n_5657_o_0),
    .Y(n_5943_o_0));
 OAI21xp33_ASAP7_75t_R n_5944 (.A1(n_5911_o_0),
    .A2(n_5923_o_0),
    .B(n_5943_o_0),
    .Y(n_5944_o_0));
 OAI21xp33_ASAP7_75t_R n_5945 (.A1(n_5790_o_0),
    .A2(n_5618_o_0),
    .B(n_5524_o_0),
    .Y(n_5945_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5946 (.A1(n_5484_o_0),
    .A2(net10),
    .B(n_5549_o_0),
    .C(n_5526_o_0),
    .Y(n_5946_o_0));
 NOR2xp33_ASAP7_75t_R n_5947 (.A(n_5484_o_0),
    .B(n_5572_o_0),
    .Y(n_5947_o_0));
 AO21x1_ASAP7_75t_R n_5948 (.A1(n_5459_o_0),
    .A2(net54),
    .B(n_5776_o_0),
    .Y(n_5948_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5949 (.A1(n_5947_o_0),
    .A2(n_5948_o_0),
    .B(n_5514_o_0),
    .C(n_5558_o_0),
    .Y(n_5949_o_0));
 OAI21xp33_ASAP7_75t_R n_5950 (.A1(n_5660_o_0),
    .A2(n_5630_o_0),
    .B(n_5949_o_0),
    .Y(n_5950_o_0));
 OAI211xp5_ASAP7_75t_R n_5951 (.A1(n_5945_o_0),
    .A2(n_5946_o_0),
    .B(n_5950_o_0),
    .C(n_5510_o_0),
    .Y(n_5951_o_0));
 INVx1_ASAP7_75t_R n_5952 (.A(n_5605_o_0),
    .Y(n_5952_o_0));
 OAI211xp5_ASAP7_75t_R n_5953 (.A1(n_5514_o_0),
    .A2(n_5743_o_0),
    .B(n_5952_o_0),
    .C(n_5606_o_0),
    .Y(n_5953_o_0));
 AOI21xp33_ASAP7_75t_R n_5954 (.A1(n_5743_o_0),
    .A2(n_5668_o_0),
    .B(n_5557_o_0),
    .Y(n_5954_o_0));
 OAI21xp33_ASAP7_75t_R n_5955 (.A1(n_5609_o_0),
    .A2(n_5501_o_0),
    .B(n_5954_o_0),
    .Y(n_5955_o_0));
 NAND3xp33_ASAP7_75t_R n_5956 (.A(n_5953_o_0),
    .B(n_5955_o_0),
    .C(n_5555_o_0),
    .Y(n_5956_o_0));
 OAI21xp33_ASAP7_75t_R n_5957 (.A1(n_5666_o_0),
    .A2(n_5577_o_0),
    .B(n_5571_o_0),
    .Y(n_5957_o_0));
 OAI311xp33_ASAP7_75t_R n_5958 (.A1(net7),
    .A2(n_5514_o_0),
    .A3(n_5549_o_0),
    .B1(n_5523_o_0),
    .C1(n_5957_o_0),
    .Y(n_5958_o_0));
 AOI31xp33_ASAP7_75t_R n_5959 (.A1(n_5514_o_0),
    .A2(n_5551_o_0),
    .A3(n_5490_o_0),
    .B(n_5523_o_0),
    .Y(n_5959_o_0));
 OAI21xp33_ASAP7_75t_R n_5960 (.A1(n_5660_o_0),
    .A2(n_5666_o_0),
    .B(n_5959_o_0),
    .Y(n_5960_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5961 (.A1(n_5571_o_0),
    .A2(n_5737_o_0),
    .B(n_5952_o_0),
    .C(n_5534_o_0),
    .Y(n_5961_o_0));
 OAI311xp33_ASAP7_75t_R n_5962 (.A1(n_5526_o_0),
    .A2(n_5685_o_0),
    .A3(n_5543_o_0),
    .B1(n_5651_o_0),
    .C1(n_5524_o_0),
    .Y(n_5962_o_0));
 AOI321xp33_ASAP7_75t_R n_5963 (.A1(n_5555_o_0),
    .A2(n_5958_o_0),
    .A3(n_5960_o_0),
    .B1(n_5961_o_0),
    .B2(n_5962_o_0),
    .C(n_5602_o_0),
    .Y(n_5963_o_0));
 AOI31xp33_ASAP7_75t_R n_5964 (.A1(n_5568_o_0),
    .A2(n_5951_o_0),
    .A3(n_5956_o_0),
    .B(n_5963_o_0),
    .Y(n_5964_o_0));
 OAI22xp33_ASAP7_75t_R n_5965 (.A1(n_5828_o_0),
    .A2(n_5571_o_0),
    .B1(n_5526_o_0),
    .B2(n_5484_o_0),
    .Y(n_5965_o_0));
 NOR3xp33_ASAP7_75t_R n_5966 (.A(n_5658_o_0),
    .B(n_5550_o_0),
    .C(n_5526_o_0),
    .Y(n_5966_o_0));
 OAI21xp33_ASAP7_75t_R n_5967 (.A1(n_5719_o_0),
    .A2(n_5966_o_0),
    .B(n_5557_o_0),
    .Y(n_5967_o_0));
 OA21x2_ASAP7_75t_R n_5968 (.A1(n_5523_o_0),
    .A2(n_5965_o_0),
    .B(n_5967_o_0),
    .Y(n_5968_o_0));
 AOI21xp33_ASAP7_75t_R n_5969 (.A1(n_5659_o_0),
    .A2(n_5591_o_0),
    .B(n_5684_o_0),
    .Y(n_5969_o_0));
 OAI21xp33_ASAP7_75t_R n_5970 (.A1(n_5571_o_0),
    .A2(n_5610_o_0),
    .B(n_5524_o_0),
    .Y(n_5970_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_5971 (.A1(n_5459_o_0),
    .A2(n_5578_o_0),
    .B(n_5597_o_0),
    .C(n_5970_o_0),
    .Y(n_5971_o_0));
 AOI21xp33_ASAP7_75t_R n_5972 (.A1(n_5557_o_0),
    .A2(n_5969_o_0),
    .B(n_5971_o_0),
    .Y(n_5972_o_0));
 OAI21xp33_ASAP7_75t_R n_5973 (.A1(n_5589_o_0),
    .A2(n_5972_o_0),
    .B(n_5567_o_0),
    .Y(n_5973_o_0));
 INVx1_ASAP7_75t_R n_5974 (.A(n_5606_o_0),
    .Y(n_5974_o_0));
 NAND3xp33_ASAP7_75t_R n_5975 (.A(n_5551_o_0),
    .B(n_5514_o_0),
    .C(n_5483_o_0),
    .Y(n_5975_o_0));
 OAI31xp33_ASAP7_75t_R n_5976 (.A1(n_5974_o_0),
    .A2(n_5744_o_0),
    .A3(n_5502_o_0),
    .B(n_5975_o_0),
    .Y(n_5976_o_0));
 OAI21xp33_ASAP7_75t_R n_5977 (.A1(n_5939_o_0),
    .A2(n_5826_o_0),
    .B(n_5844_o_0),
    .Y(n_5977_o_0));
 AOI21xp33_ASAP7_75t_R n_5978 (.A1(n_5557_o_0),
    .A2(n_5977_o_0),
    .B(n_5555_o_0),
    .Y(n_5978_o_0));
 OAI21xp33_ASAP7_75t_R n_5979 (.A1(n_5523_o_0),
    .A2(n_5976_o_0),
    .B(n_5978_o_0),
    .Y(n_5979_o_0));
 AOI21xp33_ASAP7_75t_R n_5980 (.A1(net54),
    .A2(n_5576_o_0),
    .B(n_5844_o_0),
    .Y(n_5980_o_0));
 AOI31xp33_ASAP7_75t_R n_5981 (.A1(n_5501_o_0),
    .A2(n_5547_o_0),
    .A3(n_5743_o_0),
    .B(n_5980_o_0),
    .Y(n_5981_o_0));
 OAI221xp5_ASAP7_75t_R n_5982 (.A1(n_5484_o_0),
    .A2(n_5622_o_0),
    .B1(net54),
    .B2(n_5581_o_0),
    .C(n_5571_o_0),
    .Y(n_5982_o_0));
 OAI31xp33_ASAP7_75t_R n_5983 (.A1(n_5571_o_0),
    .A2(n_5554_o_0),
    .A3(n_5666_o_0),
    .B(n_5982_o_0),
    .Y(n_5983_o_0));
 AOI21xp33_ASAP7_75t_R n_5984 (.A1(n_5558_o_0),
    .A2(n_5983_o_0),
    .B(n_5510_o_0),
    .Y(n_5984_o_0));
 OAI21xp33_ASAP7_75t_R n_5985 (.A1(n_5524_o_0),
    .A2(n_5981_o_0),
    .B(n_5984_o_0),
    .Y(n_5985_o_0));
 AOI31xp33_ASAP7_75t_R n_5986 (.A1(n_5602_o_0),
    .A2(n_5979_o_0),
    .A3(n_5985_o_0),
    .B(n_5645_o_0),
    .Y(n_5986_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_5987 (.A1(n_5968_o_0),
    .A2(n_5510_o_0),
    .B(n_5973_o_0),
    .C(n_5986_o_0),
    .Y(n_5987_o_0));
 OA21x2_ASAP7_75t_R n_5988 (.A1(n_5443_o_0),
    .A2(n_5964_o_0),
    .B(n_5987_o_0),
    .Y(n_5988_o_0));
 XNOR2xp5_ASAP7_75t_R n_5989 (.A(_01088_),
    .B(_01089_),
    .Y(n_5989_o_0));
 XNOR2xp5_ASAP7_75t_R n_5990 (.A(_01097_),
    .B(n_5989_o_0),
    .Y(n_5990_o_0));
 XOR2xp5_ASAP7_75t_R n_5991 (.A(_01010_),
    .B(_01049_),
    .Y(n_5991_o_0));
 NOR2xp33_ASAP7_75t_R n_5992 (.A(n_5991_o_0),
    .B(n_5990_o_0),
    .Y(n_5992_o_0));
 NOR2xp33_ASAP7_75t_R n_5993 (.A(_00675_),
    .B(net),
    .Y(n_5993_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_5994 (.A1(n_5990_o_0),
    .A2(n_5991_o_0),
    .B(n_5992_o_0),
    .C(net),
    .D(n_5993_o_0),
    .Y(n_5994_o_0));
 XNOR2xp5_ASAP7_75t_R n_5995 (.A(_00914_),
    .B(n_5994_o_0),
    .Y(n_5995_o_0));
 XNOR2xp5_ASAP7_75t_R n_5996 (.A(_01086_),
    .B(_01090_),
    .Y(n_5996_o_0));
 XOR2xp5_ASAP7_75t_R n_5997 (.A(n_3691_o_0),
    .B(n_5996_o_0),
    .Y(n_5997_o_0));
 XNOR2xp5_ASAP7_75t_R n_5998 (.A(_01008_),
    .B(n_3690_o_0),
    .Y(n_5998_o_0));
 NOR2xp33_ASAP7_75t_R n_5999 (.A(n_5998_o_0),
    .B(n_5997_o_0),
    .Y(n_5999_o_0));
 NOR2xp33_ASAP7_75t_R n_6000 (.A(_00677_),
    .B(net),
    .Y(n_6000_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6001 (.A1(n_5997_o_0),
    .A2(n_5998_o_0),
    .B(n_5999_o_0),
    .C(net),
    .D(n_6000_o_0),
    .Y(n_6001_o_0));
 XNOR2xp5_ASAP7_75t_R n_6002 (.A(_00912_),
    .B(n_6001_o_0),
    .Y(n_6002_o_0));
 INVx1_ASAP7_75t_R n_6003 (.A(n_6002_o_0),
    .Y(n_6003_o_0));
 XNOR2xp5_ASAP7_75t_R n_6004 (.A(_01083_),
    .B(_01090_),
    .Y(n_6004_o_0));
 INVx1_ASAP7_75t_R n_6005 (.A(n_6004_o_0),
    .Y(n_6005_o_0));
 XOR2xp5_ASAP7_75t_R n_6006 (.A(_01051_),
    .B(_01091_),
    .Y(n_6006_o_0));
 NAND2xp33_ASAP7_75t_R n_6007 (.A(n_3653_o_0),
    .B(n_6006_o_0),
    .Y(n_6007_o_0));
 OAI21xp33_ASAP7_75t_R n_6008 (.A1(n_6006_o_0),
    .A2(n_3653_o_0),
    .B(n_6007_o_0),
    .Y(n_6008_o_0));
 NOR2xp33_ASAP7_75t_R n_6009 (.A(n_3653_o_0),
    .B(n_6006_o_0),
    .Y(n_6009_o_0));
 AOI211xp5_ASAP7_75t_R n_6010 (.A1(n_6006_o_0),
    .A2(n_3653_o_0),
    .B(n_6009_o_0),
    .C(n_6005_o_0),
    .Y(n_6010_o_0));
 NOR2xp33_ASAP7_75t_R n_6011 (.A(_00540_),
    .B(net77),
    .Y(n_6011_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6012 (.A1(n_6005_o_0),
    .A2(n_6008_o_0),
    .B(n_6010_o_0),
    .C(net77),
    .D(n_6011_o_0),
    .Y(n_6012_o_0));
 OAI211xp5_ASAP7_75t_R n_6013 (.A1(n_6006_o_0),
    .A2(n_3653_o_0),
    .B(n_6007_o_0),
    .C(n_6004_o_0),
    .Y(n_6013_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6014 (.A1(n_6006_o_0),
    .A2(n_3653_o_0),
    .B(n_6009_o_0),
    .C(n_6005_o_0),
    .Y(n_6014_o_0));
 INVx1_ASAP7_75t_R n_6015 (.A(n_6011_o_0),
    .Y(n_6015_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6016 (.A1(n_6013_o_0),
    .A2(n_6014_o_0),
    .B(net3),
    .C(n_6015_o_0),
    .D(_00908_),
    .Y(n_6016_o_0));
 AO21x1_ASAP7_75t_R n_6017 (.A1(_00908_),
    .A2(n_6012_o_0),
    .B(n_6016_o_0),
    .Y(n_6017_o_0));
 XOR2xp5_ASAP7_75t_R n_6018 (.A(_01084_),
    .B(_01092_),
    .Y(n_6018_o_0));
 XNOR2xp5_ASAP7_75t_R n_6019 (.A(n_6004_o_0),
    .B(n_6018_o_0),
    .Y(n_6019_o_0));
 XNOR2xp5_ASAP7_75t_R n_6020 (.A(_01005_),
    .B(n_3647_o_0),
    .Y(n_6020_o_0));
 NAND2xp33_ASAP7_75t_R n_6021 (.A(n_6020_o_0),
    .B(n_6019_o_0),
    .Y(n_6021_o_0));
 OAI21xp33_ASAP7_75t_R n_6022 (.A1(n_6019_o_0),
    .A2(n_6020_o_0),
    .B(n_6021_o_0),
    .Y(n_6022_o_0));
 NOR2xp33_ASAP7_75t_R n_6023 (.A(_00539_),
    .B(net39),
    .Y(n_6023_o_0));
 AOI21xp33_ASAP7_75t_R n_6024 (.A1(net77),
    .A2(n_6022_o_0),
    .B(n_6023_o_0),
    .Y(n_6024_o_0));
 NOR2xp33_ASAP7_75t_R n_6025 (.A(n_6018_o_0),
    .B(n_6005_o_0),
    .Y(n_6025_o_0));
 XOR2xp5_ASAP7_75t_R n_6026 (.A(_01005_),
    .B(n_3647_o_0),
    .Y(n_6026_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6027 (.A1(n_6005_o_0),
    .A2(n_6018_o_0),
    .B(n_6025_o_0),
    .C(n_6026_o_0),
    .Y(n_6027_o_0));
 OR2x2_ASAP7_75t_R n_6028 (.A(_00539_),
    .B(net77),
    .Y(n_6028_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6029 (.A1(n_6027_o_0),
    .A2(n_6021_o_0),
    .B(net3),
    .C(n_6028_o_0),
    .D(_00909_),
    .Y(n_6029_o_0));
 AOI21x1_ASAP7_75t_R n_6030 (.A1(_00909_),
    .A2(n_6024_o_0),
    .B(n_6029_o_0),
    .Y(n_6030_o_0));
 AOI21x1_ASAP7_75t_R n_6031 (.A1(_00908_),
    .A2(n_6012_o_0),
    .B(n_6016_o_0),
    .Y(n_6031_o_0));
 INVx1_ASAP7_75t_R n_6032 (.A(_01006_),
    .Y(n_6032_o_0));
 NAND2xp33_ASAP7_75t_R n_6033 (.A(n_6032_o_0),
    .B(n_3631_o_0),
    .Y(n_6033_o_0));
 OAI21xp33_ASAP7_75t_R n_6034 (.A1(n_3631_o_0),
    .A2(n_6032_o_0),
    .B(n_6033_o_0),
    .Y(n_6034_o_0));
 NOR2xp33_ASAP7_75t_R n_6035 (.A(n_6032_o_0),
    .B(n_3631_o_0),
    .Y(n_6035_o_0));
 AOI211xp5_ASAP7_75t_R n_6036 (.A1(n_3631_o_0),
    .A2(n_6032_o_0),
    .B(n_6035_o_0),
    .C(n_3646_o_0),
    .Y(n_6036_o_0));
 NOR2xp33_ASAP7_75t_R n_6037 (.A(_00542_),
    .B(_00858_),
    .Y(n_6037_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6038 (.A1(n_3646_o_0),
    .A2(n_6034_o_0),
    .B(n_6036_o_0),
    .C(_00858_),
    .D(n_6037_o_0),
    .Y(n_6038_o_0));
 XNOR2x1_ASAP7_75t_R n_6039 (.B(n_6038_o_0),
    .Y(n_6039_o_0),
    .A(_00910_));
 NAND2xp33_ASAP7_75t_R n_6040 (.A(n_6031_o_0),
    .B(n_6039_o_0),
    .Y(n_6040_o_0));
 INVx1_ASAP7_75t_R n_6041 (.A(n_6040_o_0),
    .Y(n_6041_o_0));
 XNOR2xp5_ASAP7_75t_R n_6042 (.A(_01085_),
    .B(_01090_),
    .Y(n_6042_o_0));
 XNOR2xp5_ASAP7_75t_R n_6043 (.A(n_3617_o_0),
    .B(n_6042_o_0),
    .Y(n_6043_o_0));
 XOR2xp5_ASAP7_75t_R n_6044 (.A(_01007_),
    .B(n_3616_o_0),
    .Y(n_6044_o_0));
 NAND2xp33_ASAP7_75t_R n_6045 (.A(n_6043_o_0),
    .B(n_6044_o_0),
    .Y(n_6045_o_0));
 OAI21xp33_ASAP7_75t_R n_6046 (.A1(n_6043_o_0),
    .A2(n_6044_o_0),
    .B(n_6045_o_0),
    .Y(n_6046_o_0));
 NOR2xp33_ASAP7_75t_R n_6047 (.A(_00678_),
    .B(_00858_),
    .Y(n_6047_o_0));
 AO21x1_ASAP7_75t_R n_6048 (.A1(n_6046_o_0),
    .A2(net),
    .B(n_6047_o_0),
    .Y(n_6048_o_0));
 AOI211xp5_ASAP7_75t_R n_6049 (.A1(n_6046_o_0),
    .A2(net77),
    .B(_00911_),
    .C(n_6047_o_0),
    .Y(n_6049_o_0));
 AOI21xp5_ASAP7_75t_R n_6050 (.A1(_00911_),
    .A2(n_6048_o_0),
    .B(n_6049_o_0),
    .Y(n_6050_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6051 (.A1(n_6017_o_0),
    .A2(n_6030_o_0),
    .B(n_6041_o_0),
    .C(n_6050_o_0),
    .Y(n_6051_o_0));
 NAND2xp33_ASAP7_75t_R n_6052 (.A(n_6017_o_0),
    .B(n_6030_o_0),
    .Y(n_6052_o_0));
 NAND2xp33_ASAP7_75t_R n_6053 (.A(n_6031_o_0),
    .B(n_6039_o_0),
    .Y(n_6053_o_0));
 AOI211xp5_ASAP7_75t_R n_6054 (.A1(n_6046_o_0),
    .A2(net39),
    .B(n_868_o_0),
    .C(n_6047_o_0),
    .Y(n_6054_o_0));
 AOI21x1_ASAP7_75t_R n_6055 (.A1(n_868_o_0),
    .A2(n_6048_o_0),
    .B(n_6054_o_0),
    .Y(n_6055_o_0));
 NAND3xp33_ASAP7_75t_R n_6056 (.A(n_6052_o_0),
    .B(n_6053_o_0),
    .C(n_6055_o_0),
    .Y(n_6056_o_0));
 NAND3xp33_ASAP7_75t_R n_6057 (.A(n_6030_o_0),
    .B(n_6039_o_0),
    .C(n_6031_o_0),
    .Y(n_6057_o_0));
 XOR2x1_ASAP7_75t_R n_6058 (.A(_00910_),
    .Y(n_6058_o_0),
    .B(n_6038_o_0));
 NOR2xp33_ASAP7_75t_R n_6059 (.A(n_6020_o_0),
    .B(n_6019_o_0),
    .Y(n_6059_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6060 (.A1(n_6019_o_0),
    .A2(n_6020_o_0),
    .B(n_6059_o_0),
    .C(net),
    .Y(n_6060_o_0));
 OAI211xp5_ASAP7_75t_R n_6061 (.A1(_00539_),
    .A2(net),
    .B(n_6060_o_0),
    .C(_00909_),
    .Y(n_6061_o_0));
 OAI21xp5_ASAP7_75t_R n_6062 (.A1(_00909_),
    .A2(n_6024_o_0),
    .B(n_6061_o_0),
    .Y(n_6062_o_0));
 AOI211xp5_ASAP7_75t_R n_6063 (.A1(n_6022_o_0),
    .A2(net),
    .B(n_853_o_0),
    .C(n_6023_o_0),
    .Y(n_6063_o_0));
 OAI21xp33_ASAP7_75t_R n_6064 (.A1(n_6029_o_0),
    .A2(n_6063_o_0),
    .B(n_6017_o_0),
    .Y(n_6064_o_0));
 OAI21xp33_ASAP7_75t_R n_6065 (.A1(n_6017_o_0),
    .A2(n_6062_o_0),
    .B(n_6064_o_0),
    .Y(n_6065_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6066 (.A1(n_6046_o_0),
    .A2(net),
    .B(n_6047_o_0),
    .C(_00911_),
    .Y(n_6066_o_0));
 OAI21xp5_ASAP7_75t_R n_6067 (.A1(_00911_),
    .A2(n_6048_o_0),
    .B(n_6066_o_0),
    .Y(n_6067_o_0));
 AOI21xp33_ASAP7_75t_R n_6068 (.A1(n_6058_o_0),
    .A2(n_6065_o_0),
    .B(n_6067_o_0),
    .Y(n_6068_o_0));
 INVx1_ASAP7_75t_R n_6069 (.A(n_6029_o_0),
    .Y(n_6069_o_0));
 AOI211xp5_ASAP7_75t_R n_6070 (.A1(n_6069_o_0),
    .A2(n_6061_o_0),
    .B(n_6017_o_0),
    .C(n_6039_o_0),
    .Y(n_6070_o_0));
 OAI21xp33_ASAP7_75t_R n_6071 (.A1(n_6029_o_0),
    .A2(n_6063_o_0),
    .B(n_6017_o_0),
    .Y(n_6071_o_0));
 NOR2xp33_ASAP7_75t_R n_6072 (.A(n_6058_o_0),
    .B(n_6071_o_0),
    .Y(n_6072_o_0));
 NOR2xp33_ASAP7_75t_R n_6073 (.A(n_6070_o_0),
    .B(n_6072_o_0),
    .Y(n_6073_o_0));
 NAND2xp33_ASAP7_75t_R n_6074 (.A(_00912_),
    .B(n_6001_o_0),
    .Y(n_6074_o_0));
 OA21x2_ASAP7_75t_R n_6075 (.A1(_00912_),
    .A2(n_6001_o_0),
    .B(n_6074_o_0),
    .Y(n_6075_o_0));
 AOI221xp5_ASAP7_75t_R n_6076 (.A1(n_6057_o_0),
    .A2(n_6068_o_0),
    .B1(n_6055_o_0),
    .B2(n_6073_o_0),
    .C(n_6075_o_0),
    .Y(n_6076_o_0));
 AOI31xp33_ASAP7_75t_R n_6077 (.A1(n_6003_o_0),
    .A2(n_6051_o_0),
    .A3(n_6056_o_0),
    .B(n_6076_o_0),
    .Y(n_6077_o_0));
 AOI211xp5_ASAP7_75t_R n_6078 (.A1(n_6024_o_0),
    .A2(_00909_),
    .B(n_6031_o_0),
    .C(n_6029_o_0),
    .Y(n_6078_o_0));
 OAI21xp33_ASAP7_75t_R n_6079 (.A1(n_6039_o_0),
    .A2(n_6078_o_0),
    .B(n_6055_o_0),
    .Y(n_6079_o_0));
 INVx1_ASAP7_75t_R n_6080 (.A(n_6079_o_0),
    .Y(n_6080_o_0));
 OAI21xp33_ASAP7_75t_R n_6081 (.A1(n_6052_o_0),
    .A2(n_6058_o_0),
    .B(n_6080_o_0),
    .Y(n_6081_o_0));
 OAI21xp33_ASAP7_75t_R n_6082 (.A1(n_6058_o_0),
    .A2(n_6031_o_0),
    .B(n_6050_o_0),
    .Y(n_6082_o_0));
 AO21x1_ASAP7_75t_R n_6083 (.A1(n_6081_o_0),
    .A2(n_6082_o_0),
    .B(n_6003_o_0),
    .Y(n_6083_o_0));
 NAND3xp33_ASAP7_75t_R n_6084 (.A(n_6030_o_0),
    .B(n_6017_o_0),
    .C(n_6039_o_0),
    .Y(n_6084_o_0));
 INVx1_ASAP7_75t_R n_6085 (.A(n_6084_o_0),
    .Y(n_6085_o_0));
 NOR2xp67_ASAP7_75t_R n_6086 (.A(n_6031_o_0),
    .B(n_6039_o_0),
    .Y(n_6086_o_0));
 OAI211xp5_ASAP7_75t_R n_6087 (.A1(_00909_),
    .A2(n_6024_o_0),
    .B(n_6061_o_0),
    .C(n_6031_o_0),
    .Y(n_6087_o_0));
 AOI21xp33_ASAP7_75t_R n_6088 (.A1(n_6064_o_0),
    .A2(n_6087_o_0),
    .B(n_6039_o_0),
    .Y(n_6088_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6089 (.A1(n_6030_o_0),
    .A2(n_6031_o_0),
    .B(n_6058_o_0),
    .C(n_6055_o_0),
    .Y(n_6089_o_0));
 OAI22xp33_ASAP7_75t_R n_6090 (.A1(n_6085_o_0),
    .A2(n_6086_o_0),
    .B1(n_6088_o_0),
    .B2(n_6089_o_0),
    .Y(n_6090_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6091 (.A1(n_6046_o_0),
    .A2(net),
    .B(n_6047_o_0),
    .C(n_868_o_0),
    .Y(n_6091_o_0));
 OAI21xp5_ASAP7_75t_R n_6092 (.A1(n_868_o_0),
    .A2(n_6048_o_0),
    .B(n_6091_o_0),
    .Y(n_6092_o_0));
 NOR3xp33_ASAP7_75t_R n_6093 (.A(n_6088_o_0),
    .B(n_6092_o_0),
    .C(n_6089_o_0),
    .Y(n_6093_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6094 (.A1(n_6090_o_0),
    .A2(n_6092_o_0),
    .B(n_6093_o_0),
    .C(n_6003_o_0),
    .Y(n_6094_o_0));
 NAND2xp33_ASAP7_75t_R n_6095 (.A(_00914_),
    .B(n_5994_o_0),
    .Y(n_6095_o_0));
 OAI21xp33_ASAP7_75t_R n_6096 (.A1(_00914_),
    .A2(n_5994_o_0),
    .B(n_6095_o_0),
    .Y(n_6096_o_0));
 XNOR2xp5_ASAP7_75t_R n_6097 (.A(_01089_),
    .B(_01090_),
    .Y(n_6097_o_0));
 XNOR2xp5_ASAP7_75t_R n_6098 (.A(_01098_),
    .B(n_6097_o_0),
    .Y(n_6098_o_0));
 XOR2xp5_ASAP7_75t_R n_6099 (.A(_01011_),
    .B(_01050_),
    .Y(n_6099_o_0));
 NOR2xp33_ASAP7_75t_R n_6100 (.A(n_6099_o_0),
    .B(n_6098_o_0),
    .Y(n_6100_o_0));
 NOR2xp33_ASAP7_75t_R n_6101 (.A(_00674_),
    .B(net),
    .Y(n_6101_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6102 (.A1(n_6098_o_0),
    .A2(n_6099_o_0),
    .B(n_6100_o_0),
    .C(net),
    .D(n_6101_o_0),
    .Y(n_6102_o_0));
 NOR2xp33_ASAP7_75t_R n_6103 (.A(_00915_),
    .B(n_6102_o_0),
    .Y(n_6103_o_0));
 AOI21xp33_ASAP7_75t_R n_6104 (.A1(_00915_),
    .A2(n_6102_o_0),
    .B(n_6103_o_0),
    .Y(n_6104_o_0));
 INVx1_ASAP7_75t_R n_6105 (.A(n_6104_o_0),
    .Y(n_6105_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6106 (.A1(n_6083_o_0),
    .A2(n_6094_o_0),
    .B(n_6096_o_0),
    .C(n_6105_o_0),
    .Y(n_6106_o_0));
 INVx1_ASAP7_75t_R n_6107 (.A(n_5995_o_0),
    .Y(n_6107_o_0));
 AOI21xp33_ASAP7_75t_R n_6108 (.A1(n_6058_o_0),
    .A2(n_6030_o_0),
    .B(n_6050_o_0),
    .Y(n_6108_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6109 (.A1(n_6029_o_0),
    .A2(n_6063_o_0),
    .B(n_6031_o_0),
    .C(n_6058_o_0),
    .Y(n_6109_o_0));
 INVx1_ASAP7_75t_R n_6110 (.A(n_6109_o_0),
    .Y(n_6110_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6111 (.A1(n_6067_o_0),
    .A2(n_6031_o_0),
    .B(n_6108_o_0),
    .C(n_6110_o_0),
    .Y(n_6111_o_0));
 INVx1_ASAP7_75t_R n_6112 (.A(n_6111_o_0),
    .Y(n_6112_o_0));
 NOR3xp33_ASAP7_75t_R n_6113 (.A(n_6067_o_0),
    .B(n_6071_o_0),
    .C(n_6039_o_0),
    .Y(n_6113_o_0));
 OAI21xp33_ASAP7_75t_R n_6114 (.A1(n_6029_o_0),
    .A2(n_6063_o_0),
    .B(n_6031_o_0),
    .Y(n_6114_o_0));
 OAI21xp33_ASAP7_75t_R n_6115 (.A1(n_6058_o_0),
    .A2(n_6114_o_0),
    .B(n_6092_o_0),
    .Y(n_6115_o_0));
 OAI31xp33_ASAP7_75t_R n_6116 (.A1(n_6071_o_0),
    .A2(n_6050_o_0),
    .A3(n_6039_o_0),
    .B(n_6075_o_0),
    .Y(n_6116_o_0));
 INVx1_ASAP7_75t_R n_6117 (.A(n_6116_o_0),
    .Y(n_6117_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6118 (.A1(n_6030_o_0),
    .A2(n_6086_o_0),
    .B(n_6115_o_0),
    .C(n_6117_o_0),
    .Y(n_6118_o_0));
 OAI31xp33_ASAP7_75t_R n_6119 (.A1(n_6075_o_0),
    .A2(n_6112_o_0),
    .A3(n_6113_o_0),
    .B(n_6118_o_0),
    .Y(n_6119_o_0));
 NOR2xp33_ASAP7_75t_R n_6120 (.A(n_6058_o_0),
    .B(n_6114_o_0),
    .Y(n_6120_o_0));
 OAI31xp33_ASAP7_75t_R n_6121 (.A1(n_6050_o_0),
    .A2(n_6120_o_0),
    .A3(n_6086_o_0),
    .B(n_6002_o_0),
    .Y(n_6121_o_0));
 AOI21xp33_ASAP7_75t_R n_6122 (.A1(n_6061_o_0),
    .A2(n_6069_o_0),
    .B(n_6031_o_0),
    .Y(n_6122_o_0));
 AOI211xp5_ASAP7_75t_R n_6123 (.A1(n_6024_o_0),
    .A2(_00909_),
    .B(n_6017_o_0),
    .C(n_6029_o_0),
    .Y(n_6123_o_0));
 NOR3xp33_ASAP7_75t_R n_6124 (.A(n_6122_o_0),
    .B(n_6123_o_0),
    .C(n_6058_o_0),
    .Y(n_6124_o_0));
 OAI21xp33_ASAP7_75t_R n_6125 (.A1(n_6039_o_0),
    .A2(n_6062_o_0),
    .B(n_6092_o_0),
    .Y(n_6125_o_0));
 NOR2xp33_ASAP7_75t_R n_6126 (.A(n_6124_o_0),
    .B(n_6125_o_0),
    .Y(n_6126_o_0));
 AOI21xp33_ASAP7_75t_R n_6127 (.A1(n_6017_o_0),
    .A2(n_6062_o_0),
    .B(n_6058_o_0),
    .Y(n_6127_o_0));
 OAI21xp33_ASAP7_75t_R n_6128 (.A1(n_6127_o_0),
    .A2(n_6113_o_0),
    .B(n_6050_o_0),
    .Y(n_6128_o_0));
 AOI31xp33_ASAP7_75t_R n_6129 (.A1(n_6003_o_0),
    .A2(n_6128_o_0),
    .A3(n_6079_o_0),
    .B(n_6096_o_0),
    .Y(n_6129_o_0));
 INVx1_ASAP7_75t_R n_6130 (.A(_00915_),
    .Y(n_6130_o_0));
 NAND2xp33_ASAP7_75t_R n_6131 (.A(n_6130_o_0),
    .B(n_6102_o_0),
    .Y(n_6131_o_0));
 OAI21xp33_ASAP7_75t_R n_6132 (.A1(n_6102_o_0),
    .A2(n_6130_o_0),
    .B(n_6131_o_0),
    .Y(n_6132_o_0));
 INVx1_ASAP7_75t_R n_6133 (.A(n_6132_o_0),
    .Y(n_6133_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6134 (.A1(n_6121_o_0),
    .A2(n_6126_o_0),
    .B(n_6129_o_0),
    .C(n_6133_o_0),
    .Y(n_6134_o_0));
 OAI21xp33_ASAP7_75t_R n_6135 (.A1(n_6107_o_0),
    .A2(n_6119_o_0),
    .B(n_6134_o_0),
    .Y(n_6135_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6136 (.A1(n_5995_o_0),
    .A2(n_6077_o_0),
    .B(n_6106_o_0),
    .C(n_6135_o_0),
    .Y(n_6136_o_0));
 XNOR2xp5_ASAP7_75t_R n_6137 (.A(_01009_),
    .B(_01048_),
    .Y(n_6137_o_0));
 XNOR2xp5_ASAP7_75t_R n_6138 (.A(_01087_),
    .B(n_6137_o_0),
    .Y(n_6138_o_0));
 XOR2xp5_ASAP7_75t_R n_6139 (.A(n_3598_o_0),
    .B(n_6138_o_0),
    .Y(n_6139_o_0));
 NOR2xp33_ASAP7_75t_R n_6140 (.A(_00676_),
    .B(net),
    .Y(n_6140_o_0));
 AOI21xp33_ASAP7_75t_R n_6141 (.A1(net),
    .A2(n_6139_o_0),
    .B(n_6140_o_0),
    .Y(n_6141_o_0));
 XNOR2xp5_ASAP7_75t_R n_6142 (.A(_00913_),
    .B(n_6141_o_0),
    .Y(n_6142_o_0));
 NOR2xp33_ASAP7_75t_R n_6143 (.A(n_6031_o_0),
    .B(n_6039_o_0),
    .Y(n_6143_o_0));
 AOI21xp33_ASAP7_75t_R n_6144 (.A1(n_6030_o_0),
    .A2(n_6143_o_0),
    .B(n_6067_o_0),
    .Y(n_6144_o_0));
 OAI21xp33_ASAP7_75t_R n_6145 (.A1(n_6058_o_0),
    .A2(n_6078_o_0),
    .B(n_6144_o_0),
    .Y(n_6145_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6146 (.A1(n_6071_o_0),
    .A2(n_6058_o_0),
    .B(n_6041_o_0),
    .C(n_6055_o_0),
    .Y(n_6146_o_0));
 INVx1_ASAP7_75t_R n_6147 (.A(n_6071_o_0),
    .Y(n_6147_o_0));
 AOI31xp33_ASAP7_75t_R n_6148 (.A1(n_6050_o_0),
    .A2(n_6147_o_0),
    .A3(n_6039_o_0),
    .B(n_6075_o_0),
    .Y(n_6148_o_0));
 AOI321xp33_ASAP7_75t_R n_6149 (.A1(n_6058_o_0),
    .A2(n_6055_o_0),
    .A3(n_6030_o_0),
    .B1(n_6124_o_0),
    .B2(n_6050_o_0),
    .C(n_6002_o_0),
    .Y(n_6149_o_0));
 AOI31xp33_ASAP7_75t_R n_6150 (.A1(n_6145_o_0),
    .A2(n_6146_o_0),
    .A3(n_6148_o_0),
    .B(n_6149_o_0),
    .Y(n_6150_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6151 (.A1(n_6087_o_0),
    .A2(n_6064_o_0),
    .B(n_6039_o_0),
    .C(n_6055_o_0),
    .Y(n_6151_o_0));
 INVx1_ASAP7_75t_R n_6152 (.A(n_6151_o_0),
    .Y(n_6152_o_0));
 NAND2xp33_ASAP7_75t_R n_6153 (.A(n_6058_o_0),
    .B(n_6071_o_0),
    .Y(n_6153_o_0));
 AOI21xp33_ASAP7_75t_R n_6154 (.A1(n_6153_o_0),
    .A2(n_6110_o_0),
    .B(n_6067_o_0),
    .Y(n_6154_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6155 (.A1(n_6071_o_0),
    .A2(n_6058_o_0),
    .B(n_6152_o_0),
    .C(n_6154_o_0),
    .Y(n_6155_o_0));
 NAND2xp33_ASAP7_75t_R n_6156 (.A(n_6039_o_0),
    .B(n_6030_o_0),
    .Y(n_6156_o_0));
 AOI31xp33_ASAP7_75t_R n_6157 (.A1(n_6058_o_0),
    .A2(n_6087_o_0),
    .A3(n_6064_o_0),
    .B(n_6055_o_0),
    .Y(n_6157_o_0));
 OR2x2_ASAP7_75t_R n_6158 (.A(_00912_),
    .B(n_6001_o_0),
    .Y(n_6158_o_0));
 NAND2xp5_ASAP7_75t_R n_6159 (.A(n_6074_o_0),
    .B(n_6158_o_0),
    .Y(n_6159_o_0));
 AOI21xp33_ASAP7_75t_R n_6160 (.A1(n_6156_o_0),
    .A2(n_6157_o_0),
    .B(n_6159_o_0),
    .Y(n_6160_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6161 (.A1(n_6065_o_0),
    .A2(n_6039_o_0),
    .B(n_6050_o_0),
    .C(n_6160_o_0),
    .D(n_6104_o_0),
    .Y(n_6161_o_0));
 OAI21xp33_ASAP7_75t_R n_6162 (.A1(n_6003_o_0),
    .A2(n_6155_o_0),
    .B(n_6161_o_0),
    .Y(n_6162_o_0));
 OA21x2_ASAP7_75t_R n_6163 (.A1(n_6150_o_0),
    .A2(n_6133_o_0),
    .B(n_6162_o_0),
    .Y(n_6163_o_0));
 NOR2xp33_ASAP7_75t_R n_6164 (.A(n_6031_o_0),
    .B(n_6058_o_0),
    .Y(n_6164_o_0));
 NOR2xp33_ASAP7_75t_R n_6165 (.A(n_6050_o_0),
    .B(n_6164_o_0),
    .Y(n_6165_o_0));
 NAND3xp33_ASAP7_75t_R n_6166 (.A(n_6030_o_0),
    .B(n_6058_o_0),
    .C(n_6031_o_0),
    .Y(n_6166_o_0));
 NAND3xp33_ASAP7_75t_R n_6167 (.A(n_6165_o_0),
    .B(n_6166_o_0),
    .C(n_6159_o_0),
    .Y(n_6167_o_0));
 AOI211xp5_ASAP7_75t_R n_6168 (.A1(n_6058_o_0),
    .A2(n_6031_o_0),
    .B(n_6055_o_0),
    .C(n_6030_o_0),
    .Y(n_6168_o_0));
 AOI21xp33_ASAP7_75t_R n_6169 (.A1(n_6031_o_0),
    .A2(n_6030_o_0),
    .B(n_6039_o_0),
    .Y(n_6169_o_0));
 INVx1_ASAP7_75t_R n_6170 (.A(n_6165_o_0),
    .Y(n_6170_o_0));
 AOI21xp33_ASAP7_75t_R n_6171 (.A1(n_6030_o_0),
    .A2(n_6164_o_0),
    .B(n_6055_o_0),
    .Y(n_6171_o_0));
 NOR2xp33_ASAP7_75t_R n_6172 (.A(n_6039_o_0),
    .B(n_6030_o_0),
    .Y(n_6172_o_0));
 INVx1_ASAP7_75t_R n_6173 (.A(n_6172_o_0),
    .Y(n_6173_o_0));
 AOI21xp33_ASAP7_75t_R n_6174 (.A1(n_6171_o_0),
    .A2(n_6173_o_0),
    .B(n_6159_o_0),
    .Y(n_6174_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6175 (.A1(n_6169_o_0),
    .A2(n_6170_o_0),
    .B(n_6174_o_0),
    .C(n_6104_o_0),
    .Y(n_6175_o_0));
 NAND3xp33_ASAP7_75t_R n_6176 (.A(n_6050_o_0),
    .B(n_6078_o_0),
    .C(n_6039_o_0),
    .Y(n_6176_o_0));
 OAI211xp5_ASAP7_75t_R n_6177 (.A1(n_6031_o_0),
    .A2(n_6030_o_0),
    .B(n_6092_o_0),
    .C(n_6087_o_0),
    .Y(n_6177_o_0));
 OAI22xp33_ASAP7_75t_R n_6178 (.A1(n_6058_o_0),
    .A2(n_6092_o_0),
    .B1(n_6122_o_0),
    .B2(n_6123_o_0),
    .Y(n_6178_o_0));
 NOR3xp33_ASAP7_75t_R n_6179 (.A(n_6067_o_0),
    .B(n_6114_o_0),
    .C(n_6039_o_0),
    .Y(n_6179_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6180 (.A1(n_6177_o_0),
    .A2(n_6178_o_0),
    .B(n_6179_o_0),
    .C(n_6075_o_0),
    .Y(n_6180_o_0));
 AOI21xp33_ASAP7_75t_R n_6181 (.A1(n_6176_o_0),
    .A2(n_6180_o_0),
    .B(n_6105_o_0),
    .Y(n_6181_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6182 (.A1(n_6003_o_0),
    .A2(n_6168_o_0),
    .B(n_6175_o_0),
    .C(n_6181_o_0),
    .Y(n_6182_o_0));
 INVx1_ASAP7_75t_R n_6183 (.A(n_6096_o_0),
    .Y(n_6183_o_0));
 NAND2xp33_ASAP7_75t_R n_6184 (.A(_00913_),
    .B(n_6141_o_0),
    .Y(n_6184_o_0));
 OAI21xp33_ASAP7_75t_R n_6185 (.A1(_00913_),
    .A2(n_6141_o_0),
    .B(n_6184_o_0),
    .Y(n_6185_o_0));
 INVx1_ASAP7_75t_R n_6186 (.A(n_6185_o_0),
    .Y(n_6186_o_0));
 AOI31xp33_ASAP7_75t_R n_6187 (.A1(n_6167_o_0),
    .A2(n_6182_o_0),
    .A3(n_6183_o_0),
    .B(n_6186_o_0),
    .Y(n_6187_o_0));
 OAI21xp33_ASAP7_75t_R n_6188 (.A1(n_6107_o_0),
    .A2(n_6163_o_0),
    .B(n_6187_o_0),
    .Y(n_6188_o_0));
 OAI21xp33_ASAP7_75t_R n_6189 (.A1(n_6136_o_0),
    .A2(n_6142_o_0),
    .B(n_6188_o_0),
    .Y(n_6189_o_0));
 OAI211xp5_ASAP7_75t_R n_6190 (.A1(n_6065_o_0),
    .A2(n_6039_o_0),
    .B(n_6057_o_0),
    .C(n_6055_o_0),
    .Y(n_6190_o_0));
 INVx1_ASAP7_75t_R n_6191 (.A(n_6127_o_0),
    .Y(n_6191_o_0));
 OAI21xp33_ASAP7_75t_R n_6192 (.A1(n_6017_o_0),
    .A2(n_6062_o_0),
    .B(n_6058_o_0),
    .Y(n_6192_o_0));
 NAND2xp33_ASAP7_75t_R n_6193 (.A(n_6092_o_0),
    .B(n_6192_o_0),
    .Y(n_6193_o_0));
 INVx1_ASAP7_75t_R n_6194 (.A(n_6193_o_0),
    .Y(n_6194_o_0));
 INVx1_ASAP7_75t_R n_6195 (.A(n_6142_o_0),
    .Y(n_6195_o_0));
 AOI21xp33_ASAP7_75t_R n_6196 (.A1(n_6191_o_0),
    .A2(n_6194_o_0),
    .B(n_6195_o_0),
    .Y(n_6196_o_0));
 NAND4xp25_ASAP7_75t_R n_6197 (.A(n_6087_o_0),
    .B(n_6055_o_0),
    .C(n_6064_o_0),
    .D(n_6039_o_0),
    .Y(n_6197_o_0));
 INVx1_ASAP7_75t_R n_6198 (.A(n_6113_o_0),
    .Y(n_6198_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6199 (.A1(n_6153_o_0),
    .A2(n_6197_o_0),
    .B(n_6092_o_0),
    .C(n_6198_o_0),
    .Y(n_6199_o_0));
 AOI211xp5_ASAP7_75t_R n_6200 (.A1(n_6050_o_0),
    .A2(n_6041_o_0),
    .B(n_6199_o_0),
    .C(n_6142_o_0),
    .Y(n_6200_o_0));
 AOI21xp33_ASAP7_75t_R n_6201 (.A1(n_6190_o_0),
    .A2(n_6196_o_0),
    .B(n_6200_o_0),
    .Y(n_6201_o_0));
 NOR2xp33_ASAP7_75t_R n_6202 (.A(n_6058_o_0),
    .B(n_6030_o_0),
    .Y(n_6202_o_0));
 NOR2xp33_ASAP7_75t_R n_6203 (.A(n_6202_o_0),
    .B(n_6079_o_0),
    .Y(n_6203_o_0));
 OAI21xp33_ASAP7_75t_R n_6204 (.A1(n_6029_o_0),
    .A2(n_6063_o_0),
    .B(n_6039_o_0),
    .Y(n_6204_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6205 (.A1(n_6031_o_0),
    .A2(n_6039_o_0),
    .B(n_6204_o_0),
    .C(n_6067_o_0),
    .Y(n_6205_o_0));
 OAI21xp33_ASAP7_75t_R n_6206 (.A1(n_6031_o_0),
    .A2(n_6039_o_0),
    .B(n_6050_o_0),
    .Y(n_6206_o_0));
 AOI21xp33_ASAP7_75t_R n_6207 (.A1(n_6031_o_0),
    .A2(n_6030_o_0),
    .B(n_6039_o_0),
    .Y(n_6207_o_0));
 AOI21xp33_ASAP7_75t_R n_6208 (.A1(n_6017_o_0),
    .A2(n_6030_o_0),
    .B(n_6058_o_0),
    .Y(n_6208_o_0));
 OAI21xp33_ASAP7_75t_R n_6209 (.A1(n_6207_o_0),
    .A2(n_6208_o_0),
    .B(n_6055_o_0),
    .Y(n_6209_o_0));
 OAI211xp5_ASAP7_75t_R n_6210 (.A1(n_6206_o_0),
    .A2(n_6072_o_0),
    .B(n_6209_o_0),
    .C(n_6195_o_0),
    .Y(n_6210_o_0));
 OAI31xp33_ASAP7_75t_R n_6211 (.A1(n_6186_o_0),
    .A2(n_6203_o_0),
    .A3(n_6205_o_0),
    .B(n_6210_o_0),
    .Y(n_6211_o_0));
 OAI21xp33_ASAP7_75t_R n_6212 (.A1(n_6107_o_0),
    .A2(n_6211_o_0),
    .B(n_6105_o_0),
    .Y(n_6212_o_0));
 AOI21xp33_ASAP7_75t_R n_6213 (.A1(n_6183_o_0),
    .A2(n_6201_o_0),
    .B(n_6212_o_0),
    .Y(n_6213_o_0));
 NOR2xp33_ASAP7_75t_R n_6214 (.A(n_6039_o_0),
    .B(n_6030_o_0),
    .Y(n_6214_o_0));
 INVx1_ASAP7_75t_R n_6215 (.A(n_6214_o_0),
    .Y(n_6215_o_0));
 INVx1_ASAP7_75t_R n_6216 (.A(n_6176_o_0),
    .Y(n_6216_o_0));
 AOI21xp33_ASAP7_75t_R n_6217 (.A1(n_6067_o_0),
    .A2(n_6156_o_0),
    .B(n_6216_o_0),
    .Y(n_6217_o_0));
 AOI21xp33_ASAP7_75t_R n_6218 (.A1(n_6058_o_0),
    .A2(n_6065_o_0),
    .B(n_6050_o_0),
    .Y(n_6218_o_0));
 OAI21xp33_ASAP7_75t_R n_6219 (.A1(n_6039_o_0),
    .A2(n_6078_o_0),
    .B(n_6092_o_0),
    .Y(n_6219_o_0));
 OAI21xp33_ASAP7_75t_R n_6220 (.A1(n_6219_o_0),
    .A2(n_6041_o_0),
    .B(n_6186_o_0),
    .Y(n_6220_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6221 (.A1(n_6031_o_0),
    .A2(n_6058_o_0),
    .B(n_6218_o_0),
    .C(n_6220_o_0),
    .Y(n_6221_o_0));
 AOI31xp33_ASAP7_75t_R n_6222 (.A1(n_6215_o_0),
    .A2(n_6217_o_0),
    .A3(n_6142_o_0),
    .B(n_6221_o_0),
    .Y(n_6222_o_0));
 INVx1_ASAP7_75t_R n_6223 (.A(n_6153_o_0),
    .Y(n_6223_o_0));
 INVx1_ASAP7_75t_R n_6224 (.A(n_6078_o_0),
    .Y(n_6224_o_0));
 OAI21xp33_ASAP7_75t_R n_6225 (.A1(n_6058_o_0),
    .A2(n_6224_o_0),
    .B(n_6218_o_0),
    .Y(n_6225_o_0));
 OAI31xp33_ASAP7_75t_R n_6226 (.A1(n_6055_o_0),
    .A2(n_6041_o_0),
    .A3(n_6223_o_0),
    .B(n_6225_o_0),
    .Y(n_6226_o_0));
 INVx1_ASAP7_75t_R n_6227 (.A(n_6052_o_0),
    .Y(n_6227_o_0));
 NOR2xp33_ASAP7_75t_R n_6228 (.A(n_6039_o_0),
    .B(n_6055_o_0),
    .Y(n_6228_o_0));
 OAI21xp33_ASAP7_75t_R n_6229 (.A1(n_6089_o_0),
    .A2(n_6172_o_0),
    .B(n_6186_o_0),
    .Y(n_6229_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6230 (.A1(n_6227_o_0),
    .A2(n_6062_o_0),
    .B(n_6228_o_0),
    .C(n_6229_o_0),
    .Y(n_6230_o_0));
 AOI211xp5_ASAP7_75t_R n_6231 (.A1(n_6226_o_0),
    .A2(n_6185_o_0),
    .B(n_5995_o_0),
    .C(n_6230_o_0),
    .Y(n_6231_o_0));
 AOI211xp5_ASAP7_75t_R n_6232 (.A1(n_6096_o_0),
    .A2(n_6222_o_0),
    .B(n_6231_o_0),
    .C(n_6105_o_0),
    .Y(n_6232_o_0));
 NAND3xp33_ASAP7_75t_R n_6233 (.A(n_6050_o_0),
    .B(n_6078_o_0),
    .C(n_6058_o_0),
    .Y(n_6233_o_0));
 OAI31xp33_ASAP7_75t_R n_6234 (.A1(n_6086_o_0),
    .A2(n_6124_o_0),
    .A3(n_6055_o_0),
    .B(n_6142_o_0),
    .Y(n_6234_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6235 (.A1(n_6052_o_0),
    .A2(n_6030_o_0),
    .B(n_6086_o_0),
    .C(n_6055_o_0),
    .D(n_6234_o_0),
    .Y(n_6235_o_0));
 AOI311xp33_ASAP7_75t_R n_6236 (.A1(n_6195_o_0),
    .A2(n_6190_o_0),
    .A3(n_6233_o_0),
    .B(n_6096_o_0),
    .C(n_6235_o_0),
    .Y(n_6236_o_0));
 NOR2xp33_ASAP7_75t_R n_6237 (.A(n_6031_o_0),
    .B(n_6030_o_0),
    .Y(n_6237_o_0));
 INVx1_ASAP7_75t_R n_6238 (.A(n_6237_o_0),
    .Y(n_6238_o_0));
 INVx1_ASAP7_75t_R n_6239 (.A(n_6125_o_0),
    .Y(n_6239_o_0));
 AOI22xp33_ASAP7_75t_R n_6240 (.A1(n_6238_o_0),
    .A2(n_6239_o_0),
    .B1(n_6055_o_0),
    .B2(n_6208_o_0),
    .Y(n_6240_o_0));
 NAND2xp33_ASAP7_75t_R n_6241 (.A(n_6031_o_0),
    .B(n_6030_o_0),
    .Y(n_6241_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6242 (.A1(n_6087_o_0),
    .A2(n_6064_o_0),
    .B(n_6058_o_0),
    .C(n_6055_o_0),
    .Y(n_6242_o_0));
 AOI21xp33_ASAP7_75t_R n_6243 (.A1(n_6058_o_0),
    .A2(n_6241_o_0),
    .B(n_6242_o_0),
    .Y(n_6243_o_0));
 INVx1_ASAP7_75t_R n_6244 (.A(n_6145_o_0),
    .Y(n_6244_o_0));
 OAI31xp33_ASAP7_75t_R n_6245 (.A1(n_6243_o_0),
    .A2(n_6244_o_0),
    .A3(n_6186_o_0),
    .B(n_6096_o_0),
    .Y(n_6245_o_0));
 AOI21xp33_ASAP7_75t_R n_6246 (.A1(n_6186_o_0),
    .A2(n_6240_o_0),
    .B(n_6245_o_0),
    .Y(n_6246_o_0));
 NOR2xp33_ASAP7_75t_R n_6247 (.A(n_6058_o_0),
    .B(n_6030_o_0),
    .Y(n_6247_o_0));
 OAI211xp5_ASAP7_75t_R n_6248 (.A1(n_6058_o_0),
    .A2(n_6114_o_0),
    .B(n_6166_o_0),
    .C(n_6092_o_0),
    .Y(n_6248_o_0));
 OAI31xp33_ASAP7_75t_R n_6249 (.A1(n_6050_o_0),
    .A2(n_6186_o_0),
    .A3(n_6247_o_0),
    .B(n_6248_o_0),
    .Y(n_6249_o_0));
 AOI21xp33_ASAP7_75t_R n_6250 (.A1(n_6096_o_0),
    .A2(n_6249_o_0),
    .B(n_6132_o_0),
    .Y(n_6250_o_0));
 NOR2xp33_ASAP7_75t_R n_6251 (.A(n_6055_o_0),
    .B(n_6164_o_0),
    .Y(n_6251_o_0));
 AOI21xp33_ASAP7_75t_R n_6252 (.A1(n_6166_o_0),
    .A2(n_6251_o_0),
    .B(n_6195_o_0),
    .Y(n_6252_o_0));
 OAI21xp33_ASAP7_75t_R n_6253 (.A1(n_6050_o_0),
    .A2(n_6088_o_0),
    .B(n_6252_o_0),
    .Y(n_6253_o_0));
 NOR2xp33_ASAP7_75t_R n_6254 (.A(n_6017_o_0),
    .B(n_6039_o_0),
    .Y(n_6254_o_0));
 OAI21xp33_ASAP7_75t_R n_6255 (.A1(n_6031_o_0),
    .A2(n_6062_o_0),
    .B(n_6058_o_0),
    .Y(n_6255_o_0));
 AOI21xp33_ASAP7_75t_R n_6256 (.A1(n_6062_o_0),
    .A2(n_6039_o_0),
    .B(n_6050_o_0),
    .Y(n_6256_o_0));
 AOI21xp33_ASAP7_75t_R n_6257 (.A1(n_6255_o_0),
    .A2(n_6256_o_0),
    .B(n_6185_o_0),
    .Y(n_6257_o_0));
 OAI31xp33_ASAP7_75t_R n_6258 (.A1(n_6055_o_0),
    .A2(n_6072_o_0),
    .A3(n_6254_o_0),
    .B(n_6257_o_0),
    .Y(n_6258_o_0));
 NAND3xp33_ASAP7_75t_R n_6259 (.A(n_6253_o_0),
    .B(n_6258_o_0),
    .C(n_6107_o_0),
    .Y(n_6259_o_0));
 AOI21xp33_ASAP7_75t_R n_6260 (.A1(n_6250_o_0),
    .A2(n_6259_o_0),
    .B(n_6075_o_0),
    .Y(n_6260_o_0));
 OAI31xp33_ASAP7_75t_R n_6261 (.A1(n_6105_o_0),
    .A2(n_6236_o_0),
    .A3(n_6246_o_0),
    .B(n_6260_o_0),
    .Y(n_6261_o_0));
 OAI31xp33_ASAP7_75t_R n_6262 (.A1(n_6002_o_0),
    .A2(n_6213_o_0),
    .A3(n_6232_o_0),
    .B(n_6261_o_0),
    .Y(n_6262_o_0));
 INVx1_ASAP7_75t_R n_6263 (.A(n_6124_o_0),
    .Y(n_6263_o_0));
 NOR3xp33_ASAP7_75t_R n_6264 (.A(n_6109_o_0),
    .B(n_6086_o_0),
    .C(n_6055_o_0),
    .Y(n_6264_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6265 (.A1(n_6263_o_0),
    .A2(n_6218_o_0),
    .B(n_6264_o_0),
    .C(n_6002_o_0),
    .Y(n_6265_o_0));
 INVx1_ASAP7_75t_R n_6266 (.A(n_6204_o_0),
    .Y(n_6266_o_0));
 OAI21xp33_ASAP7_75t_R n_6267 (.A1(n_6039_o_0),
    .A2(n_6114_o_0),
    .B(n_6067_o_0),
    .Y(n_6267_o_0));
 INVx1_ASAP7_75t_R n_6268 (.A(n_6254_o_0),
    .Y(n_6268_o_0));
 AOI31xp33_ASAP7_75t_R n_6269 (.A1(n_6031_o_0),
    .A2(n_6030_o_0),
    .A3(n_6039_o_0),
    .B(n_6055_o_0),
    .Y(n_6269_o_0));
 AOI21xp33_ASAP7_75t_R n_6270 (.A1(n_6268_o_0),
    .A2(n_6269_o_0),
    .B(n_6159_o_0),
    .Y(n_6270_o_0));
 OAI21xp33_ASAP7_75t_R n_6271 (.A1(n_6266_o_0),
    .A2(n_6267_o_0),
    .B(n_6270_o_0),
    .Y(n_6271_o_0));
 NOR2xp33_ASAP7_75t_R n_6272 (.A(n_6058_o_0),
    .B(n_6078_o_0),
    .Y(n_6272_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6273 (.A1(n_6062_o_0),
    .A2(n_6092_o_0),
    .B(n_6058_o_0),
    .C(n_6272_o_0),
    .Y(n_6273_o_0));
 OAI211xp5_ASAP7_75t_R n_6274 (.A1(n_6058_o_0),
    .A2(n_6224_o_0),
    .B(n_6268_o_0),
    .C(n_6067_o_0),
    .Y(n_6274_o_0));
 OAI32xp33_ASAP7_75t_R n_6275 (.A1(n_6067_o_0),
    .A2(n_6114_o_0),
    .A3(n_6039_o_0),
    .B1(n_6269_o_0),
    .B2(n_6159_o_0),
    .Y(n_6275_o_0));
 AOI221xp5_ASAP7_75t_R n_6276 (.A1(n_6002_o_0),
    .A2(n_6273_o_0),
    .B1(n_6274_o_0),
    .B2(n_6275_o_0),
    .C(n_6186_o_0),
    .Y(n_6276_o_0));
 AOI31xp33_ASAP7_75t_R n_6277 (.A1(n_6195_o_0),
    .A2(n_6265_o_0),
    .A3(n_6271_o_0),
    .B(n_6276_o_0),
    .Y(n_6277_o_0));
 NAND2xp33_ASAP7_75t_R n_6278 (.A(n_6039_o_0),
    .B(n_6062_o_0),
    .Y(n_6278_o_0));
 OAI211xp5_ASAP7_75t_R n_6279 (.A1(n_6031_o_0),
    .A2(n_6039_o_0),
    .B(n_6278_o_0),
    .C(n_6055_o_0),
    .Y(n_6279_o_0));
 INVx1_ASAP7_75t_R n_6280 (.A(n_6279_o_0),
    .Y(n_6280_o_0));
 AOI31xp33_ASAP7_75t_R n_6281 (.A1(n_6058_o_0),
    .A2(n_6050_o_0),
    .A3(n_6030_o_0),
    .B(n_6075_o_0),
    .Y(n_6281_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6282 (.A1(n_6227_o_0),
    .A2(n_6058_o_0),
    .B(n_6242_o_0),
    .C(n_6281_o_0),
    .Y(n_6282_o_0));
 OAI31xp33_ASAP7_75t_R n_6283 (.A1(n_6280_o_0),
    .A2(n_6126_o_0),
    .A3(n_6002_o_0),
    .B(n_6282_o_0),
    .Y(n_6283_o_0));
 OAI21xp33_ASAP7_75t_R n_6284 (.A1(n_6031_o_0),
    .A2(n_6030_o_0),
    .B(n_6108_o_0),
    .Y(n_6284_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6285 (.A1(n_6055_o_0),
    .A2(n_6247_o_0),
    .B(n_6284_o_0),
    .C(n_6003_o_0),
    .Y(n_6285_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6286 (.A1(n_6123_o_0),
    .A2(n_6122_o_0),
    .B(n_6039_o_0),
    .C(n_6070_o_0),
    .Y(n_6286_o_0));
 OAI21xp33_ASAP7_75t_R n_6287 (.A1(n_6050_o_0),
    .A2(n_6286_o_0),
    .B(n_6075_o_0),
    .Y(n_6287_o_0));
 AOI21xp33_ASAP7_75t_R n_6288 (.A1(n_6239_o_0),
    .A2(n_6191_o_0),
    .B(n_6287_o_0),
    .Y(n_6288_o_0));
 OAI21xp33_ASAP7_75t_R n_6289 (.A1(n_6285_o_0),
    .A2(n_6288_o_0),
    .B(n_6142_o_0),
    .Y(n_6289_o_0));
 OAI211xp5_ASAP7_75t_R n_6290 (.A1(n_6185_o_0),
    .A2(n_6283_o_0),
    .B(n_6289_o_0),
    .C(n_6132_o_0),
    .Y(n_6290_o_0));
 OAI21xp33_ASAP7_75t_R n_6291 (.A1(n_6104_o_0),
    .A2(n_6277_o_0),
    .B(n_6290_o_0),
    .Y(n_6291_o_0));
 INVx1_ASAP7_75t_R n_6292 (.A(n_6171_o_0),
    .Y(n_6292_o_0));
 NAND3xp33_ASAP7_75t_R n_6293 (.A(n_6030_o_0),
    .B(n_6039_o_0),
    .C(n_6031_o_0),
    .Y(n_6293_o_0));
 NAND3xp33_ASAP7_75t_R n_6294 (.A(n_6192_o_0),
    .B(n_6293_o_0),
    .C(n_6067_o_0),
    .Y(n_6294_o_0));
 AOI21xp33_ASAP7_75t_R n_6295 (.A1(n_6292_o_0),
    .A2(n_6294_o_0),
    .B(n_6075_o_0),
    .Y(n_6295_o_0));
 OAI21xp33_ASAP7_75t_R n_6296 (.A1(n_6058_o_0),
    .A2(n_6071_o_0),
    .B(n_6067_o_0),
    .Y(n_6296_o_0));
 OAI21xp33_ASAP7_75t_R n_6297 (.A1(n_6254_o_0),
    .A2(n_6296_o_0),
    .B(n_6075_o_0),
    .Y(n_6297_o_0));
 AOI21xp33_ASAP7_75t_R n_6298 (.A1(n_6157_o_0),
    .A2(n_6204_o_0),
    .B(n_6297_o_0),
    .Y(n_6298_o_0));
 OAI31xp33_ASAP7_75t_R n_6299 (.A1(n_6017_o_0),
    .A2(n_6063_o_0),
    .A3(n_6029_o_0),
    .B(n_6039_o_0),
    .Y(n_6299_o_0));
 AOI321xp33_ASAP7_75t_R n_6300 (.A1(n_6092_o_0),
    .A2(n_6255_o_0),
    .A3(n_6299_o_0),
    .B1(n_6084_o_0),
    .B2(n_6108_o_0),
    .C(n_6186_o_0),
    .Y(n_6300_o_0));
 NOR2xp33_ASAP7_75t_R n_6301 (.A(n_6075_o_0),
    .B(n_6186_o_0),
    .Y(n_6301_o_0));
 NOR2xp33_ASAP7_75t_R n_6302 (.A(n_6058_o_0),
    .B(n_6078_o_0),
    .Y(n_6302_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6303 (.A1(n_6030_o_0),
    .A2(n_6086_o_0),
    .B(n_6302_o_0),
    .C(n_6055_o_0),
    .Y(n_6303_o_0));
 OAI211xp5_ASAP7_75t_R n_6304 (.A1(n_6124_o_0),
    .A2(n_6125_o_0),
    .B(n_6303_o_0),
    .C(n_6159_o_0),
    .Y(n_6304_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6305 (.A1(n_6075_o_0),
    .A2(n_6300_o_0),
    .B(n_6301_o_0),
    .C(n_6304_o_0),
    .Y(n_6305_o_0));
 OAI31xp33_ASAP7_75t_R n_6306 (.A1(n_6142_o_0),
    .A2(n_6295_o_0),
    .A3(n_6298_o_0),
    .B(n_6305_o_0),
    .Y(n_6306_o_0));
 AO21x1_ASAP7_75t_R n_6307 (.A1(n_6306_o_0),
    .A2(n_6105_o_0),
    .B(n_6107_o_0),
    .Y(n_6307_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6308 (.A1(n_6030_o_0),
    .A2(n_6058_o_0),
    .B(n_6050_o_0),
    .C(n_6292_o_0),
    .Y(n_6308_o_0));
 AOI21xp33_ASAP7_75t_R n_6309 (.A1(n_6084_o_0),
    .A2(n_6108_o_0),
    .B(n_6159_o_0),
    .Y(n_6309_o_0));
 OAI31xp33_ASAP7_75t_R n_6310 (.A1(n_6062_o_0),
    .A2(n_6058_o_0),
    .A3(n_6055_o_0),
    .B(n_6309_o_0),
    .Y(n_6310_o_0));
 OA21x2_ASAP7_75t_R n_6311 (.A1(n_6308_o_0),
    .A2(n_6003_o_0),
    .B(n_6310_o_0),
    .Y(n_6311_o_0));
 AOI21xp33_ASAP7_75t_R n_6312 (.A1(n_6058_o_0),
    .A2(n_6031_o_0),
    .B(n_6050_o_0),
    .Y(n_6312_o_0));
 INVx1_ASAP7_75t_R n_6313 (.A(n_6166_o_0),
    .Y(n_6313_o_0));
 OAI21xp33_ASAP7_75t_R n_6314 (.A1(n_6115_o_0),
    .A2(n_6313_o_0),
    .B(n_6003_o_0),
    .Y(n_6314_o_0));
 NAND3xp33_ASAP7_75t_R n_6315 (.A(n_6092_o_0),
    .B(n_6071_o_0),
    .C(n_6058_o_0),
    .Y(n_6315_o_0));
 OAI211xp5_ASAP7_75t_R n_6316 (.A1(n_6151_o_0),
    .A2(n_6272_o_0),
    .B(n_6315_o_0),
    .C(n_6159_o_0),
    .Y(n_6316_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6317 (.A1(n_6312_o_0),
    .A2(n_6057_o_0),
    .B(n_6314_o_0),
    .C(n_6316_o_0),
    .Y(n_6317_o_0));
 OAI21xp33_ASAP7_75t_R n_6318 (.A1(n_6185_o_0),
    .A2(n_6317_o_0),
    .B(n_6132_o_0),
    .Y(n_6318_o_0));
 AOI21xp33_ASAP7_75t_R n_6319 (.A1(n_6142_o_0),
    .A2(n_6311_o_0),
    .B(n_6318_o_0),
    .Y(n_6319_o_0));
 OAI22xp33_ASAP7_75t_R n_6320 (.A1(n_6291_o_0),
    .A2(n_6096_o_0),
    .B1(n_6307_o_0),
    .B2(n_6319_o_0),
    .Y(n_6320_o_0));
 INVx1_ASAP7_75t_R n_6321 (.A(n_6065_o_0),
    .Y(n_6321_o_0));
 OAI21xp33_ASAP7_75t_R n_6322 (.A1(n_6058_o_0),
    .A2(n_6114_o_0),
    .B(n_6239_o_0),
    .Y(n_6322_o_0));
 OAI31xp33_ASAP7_75t_R n_6323 (.A1(n_6050_o_0),
    .A2(n_6321_o_0),
    .A3(n_6058_o_0),
    .B(n_6322_o_0),
    .Y(n_6323_o_0));
 INVx1_ASAP7_75t_R n_6324 (.A(n_6312_o_0),
    .Y(n_6324_o_0));
 NAND2xp33_ASAP7_75t_R n_6325 (.A(n_6017_o_0),
    .B(n_6039_o_0),
    .Y(n_6325_o_0));
 NAND3xp33_ASAP7_75t_R n_6326 (.A(n_6067_o_0),
    .B(n_6087_o_0),
    .C(n_6064_o_0),
    .Y(n_6326_o_0));
 OAI22xp33_ASAP7_75t_R n_6327 (.A1(n_6058_o_0),
    .A2(n_6067_o_0),
    .B1(n_6122_o_0),
    .B2(n_6123_o_0),
    .Y(n_6327_o_0));
 AOI31xp33_ASAP7_75t_R n_6328 (.A1(n_6325_o_0),
    .A2(n_6326_o_0),
    .A3(n_6327_o_0),
    .B(n_6075_o_0),
    .Y(n_6328_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6329 (.A1(n_6039_o_0),
    .A2(n_6241_o_0),
    .B(n_6324_o_0),
    .C(n_6328_o_0),
    .Y(n_6329_o_0));
 OAI21xp33_ASAP7_75t_R n_6330 (.A1(n_6323_o_0),
    .A2(n_6116_o_0),
    .B(n_6329_o_0),
    .Y(n_6330_o_0));
 INVx1_ASAP7_75t_R n_6331 (.A(n_6114_o_0),
    .Y(n_6331_o_0));
 OAI21xp33_ASAP7_75t_R n_6332 (.A1(n_6058_o_0),
    .A2(n_6331_o_0),
    .B(n_6312_o_0),
    .Y(n_6332_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6333 (.A1(n_6115_o_0),
    .A2(n_6313_o_0),
    .B(n_6332_o_0),
    .C(n_6003_o_0),
    .Y(n_6333_o_0));
 NOR3xp33_ASAP7_75t_R n_6334 (.A(n_6333_o_0),
    .B(n_6270_o_0),
    .C(n_5995_o_0),
    .Y(n_6334_o_0));
 AOI21xp33_ASAP7_75t_R n_6335 (.A1(n_6096_o_0),
    .A2(n_6330_o_0),
    .B(n_6334_o_0),
    .Y(n_6335_o_0));
 NAND4xp25_ASAP7_75t_R n_6336 (.A(n_6055_o_0),
    .B(n_6058_o_0),
    .C(n_6062_o_0),
    .D(n_6031_o_0),
    .Y(n_6336_o_0));
 INVx1_ASAP7_75t_R n_6337 (.A(n_6336_o_0),
    .Y(n_6337_o_0));
 INVx1_ASAP7_75t_R n_6338 (.A(n_6088_o_0),
    .Y(n_6338_o_0));
 OAI21xp33_ASAP7_75t_R n_6339 (.A1(n_6067_o_0),
    .A2(n_6338_o_0),
    .B(n_6117_o_0),
    .Y(n_6339_o_0));
 OAI31xp33_ASAP7_75t_R n_6340 (.A1(n_6075_o_0),
    .A2(n_6264_o_0),
    .A3(n_6337_o_0),
    .B(n_6339_o_0),
    .Y(n_6340_o_0));
 OAI211xp5_ASAP7_75t_R n_6341 (.A1(n_6125_o_0),
    .A2(n_6237_o_0),
    .B(n_6146_o_0),
    .C(n_6159_o_0),
    .Y(n_6341_o_0));
 NAND2xp33_ASAP7_75t_R n_6342 (.A(n_6327_o_0),
    .B(n_6326_o_0),
    .Y(n_6342_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6343 (.A1(n_6058_o_0),
    .A2(n_6331_o_0),
    .B(n_6164_o_0),
    .C(n_6055_o_0),
    .D(n_6002_o_0),
    .Y(n_6343_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6344 (.A1(n_6039_o_0),
    .A2(n_6241_o_0),
    .B(n_6342_o_0),
    .C(n_6343_o_0),
    .Y(n_6344_o_0));
 AOI31xp33_ASAP7_75t_R n_6345 (.A1(n_6341_o_0),
    .A2(n_6344_o_0),
    .A3(n_6183_o_0),
    .B(n_6142_o_0),
    .Y(n_6345_o_0));
 OAI21xp33_ASAP7_75t_R n_6346 (.A1(n_6107_o_0),
    .A2(n_6340_o_0),
    .B(n_6345_o_0),
    .Y(n_6346_o_0));
 OAI21xp33_ASAP7_75t_R n_6347 (.A1(n_6186_o_0),
    .A2(n_6335_o_0),
    .B(n_6346_o_0),
    .Y(n_6347_o_0));
 OAI21xp33_ASAP7_75t_R n_6348 (.A1(n_6058_o_0),
    .A2(n_6331_o_0),
    .B(n_6068_o_0),
    .Y(n_6348_o_0));
 NAND3xp33_ASAP7_75t_R n_6349 (.A(n_6348_o_0),
    .B(n_6056_o_0),
    .C(n_6003_o_0),
    .Y(n_6349_o_0));
 AOI22xp33_ASAP7_75t_R n_6350 (.A1(n_6122_o_0),
    .A2(n_6039_o_0),
    .B1(n_6030_o_0),
    .B2(n_6031_o_0),
    .Y(n_6350_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6351 (.A1(n_6017_o_0),
    .A2(n_6039_o_0),
    .B(n_6070_o_0),
    .C(n_6256_o_0),
    .Y(n_6351_o_0));
 OAI211xp5_ASAP7_75t_R n_6352 (.A1(n_6350_o_0),
    .A2(n_6055_o_0),
    .B(n_6351_o_0),
    .C(n_6002_o_0),
    .Y(n_6352_o_0));
 OAI21xp33_ASAP7_75t_R n_6353 (.A1(n_6123_o_0),
    .A2(n_6122_o_0),
    .B(n_6039_o_0),
    .Y(n_6353_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6354 (.A1(n_6039_o_0),
    .A2(n_6114_o_0),
    .B(n_6325_o_0),
    .C(n_6055_o_0),
    .Y(n_6354_o_0));
 AOI31xp33_ASAP7_75t_R n_6355 (.A1(n_6067_o_0),
    .A2(n_6153_o_0),
    .A3(n_6353_o_0),
    .B(n_6354_o_0),
    .Y(n_6355_o_0));
 OAI311xp33_ASAP7_75t_R n_6356 (.A1(n_6039_o_0),
    .A2(n_6122_o_0),
    .A3(n_6123_o_0),
    .B1(n_6092_o_0),
    .C1(n_6204_o_0),
    .Y(n_6356_o_0));
 OAI31xp33_ASAP7_75t_R n_6357 (.A1(n_6050_o_0),
    .A2(n_6169_o_0),
    .A3(n_6302_o_0),
    .B(n_6356_o_0),
    .Y(n_6357_o_0));
 AOI321xp33_ASAP7_75t_R n_6358 (.A1(n_6158_o_0),
    .A2(n_6355_o_0),
    .A3(n_6074_o_0),
    .B1(n_6159_o_0),
    .B2(n_6357_o_0),
    .C(n_6107_o_0),
    .Y(n_6358_o_0));
 AOI31xp33_ASAP7_75t_R n_6359 (.A1(n_6107_o_0),
    .A2(n_6349_o_0),
    .A3(n_6352_o_0),
    .B(n_6358_o_0),
    .Y(n_6359_o_0));
 NAND2xp33_ASAP7_75t_R n_6360 (.A(n_6017_o_0),
    .B(n_6030_o_0),
    .Y(n_6360_o_0));
 INVx1_ASAP7_75t_R n_6361 (.A(n_6054_o_0),
    .Y(n_6361_o_0));
 AOI22xp33_ASAP7_75t_R n_6362 (.A1(n_6361_o_0),
    .A2(n_6091_o_0),
    .B1(n_6058_o_0),
    .B2(n_6031_o_0),
    .Y(n_6362_o_0));
 OAI21xp33_ASAP7_75t_R n_6363 (.A1(n_6202_o_0),
    .A2(n_6151_o_0),
    .B(n_6159_o_0),
    .Y(n_6363_o_0));
 OAI211xp5_ASAP7_75t_R n_6364 (.A1(n_6206_o_0),
    .A2(n_6202_o_0),
    .B(n_6242_o_0),
    .C(n_6003_o_0),
    .Y(n_6364_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6365 (.A1(n_6360_o_0),
    .A2(n_6362_o_0),
    .B(n_6363_o_0),
    .C(n_6364_o_0),
    .Y(n_6365_o_0));
 INVx1_ASAP7_75t_R n_6366 (.A(n_6299_o_0),
    .Y(n_6366_o_0));
 OAI311xp33_ASAP7_75t_R n_6367 (.A1(n_6039_o_0),
    .A2(n_6123_o_0),
    .A3(n_6122_o_0),
    .B1(n_6092_o_0),
    .C1(n_6110_o_0),
    .Y(n_6367_o_0));
 OAI311xp33_ASAP7_75t_R n_6368 (.A1(n_6050_o_0),
    .A2(n_6172_o_0),
    .A3(n_6366_o_0),
    .B1(n_6183_o_0),
    .C1(n_6367_o_0),
    .Y(n_6368_o_0));
 NAND2xp33_ASAP7_75t_R n_6369 (.A(n_6002_o_0),
    .B(n_6183_o_0),
    .Y(n_6369_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6370 (.A1(n_6362_o_0),
    .A2(n_6360_o_0),
    .B(n_6055_o_0),
    .C(n_6002_o_0),
    .Y(n_6370_o_0));
 AOI211xp5_ASAP7_75t_R n_6371 (.A1(n_6227_o_0),
    .A2(n_6039_o_0),
    .B(n_6370_o_0),
    .C(n_6195_o_0),
    .Y(n_6371_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6372 (.A1(n_6002_o_0),
    .A2(n_6368_o_0),
    .B(n_6369_o_0),
    .C(n_6371_o_0),
    .Y(n_6372_o_0));
 AOI311xp33_ASAP7_75t_R n_6373 (.A1(n_6058_o_0),
    .A2(n_6087_o_0),
    .A3(n_6064_o_0),
    .B(n_6055_o_0),
    .C(n_6109_o_0),
    .Y(n_6373_o_0));
 AOI31xp33_ASAP7_75t_R n_6374 (.A1(n_6067_o_0),
    .A2(n_6173_o_0),
    .A3(n_6299_o_0),
    .B(n_6373_o_0),
    .Y(n_6374_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6375 (.A1(n_6002_o_0),
    .A2(n_6374_o_0),
    .B(n_6183_o_0),
    .C(n_6142_o_0),
    .Y(n_6375_o_0));
 AOI211xp5_ASAP7_75t_R n_6376 (.A1(n_6096_o_0),
    .A2(n_6365_o_0),
    .B(n_6372_o_0),
    .C(n_6375_o_0),
    .Y(n_6376_o_0));
 AOI211xp5_ASAP7_75t_R n_6377 (.A1(n_6359_o_0),
    .A2(n_6186_o_0),
    .B(n_6376_o_0),
    .C(n_6133_o_0),
    .Y(n_6377_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6378 (.A1(_00915_),
    .A2(n_6102_o_0),
    .B(n_6103_o_0),
    .C(n_6347_o_0),
    .D(n_6377_o_0),
    .Y(n_6378_o_0));
 AOI21xp33_ASAP7_75t_R n_6379 (.A1(n_6204_o_0),
    .A2(n_6360_o_0),
    .B(n_6067_o_0),
    .Y(n_6379_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6380 (.A1(n_6109_o_0),
    .A2(n_6254_o_0),
    .B(n_6055_o_0),
    .C(n_6379_o_0),
    .Y(n_6380_o_0));
 NOR2xp33_ASAP7_75t_R n_6381 (.A(n_6109_o_0),
    .B(n_6172_o_0),
    .Y(n_6381_o_0));
 AOI22xp33_ASAP7_75t_R n_6382 (.A1(n_6381_o_0),
    .A2(n_6067_o_0),
    .B1(n_6360_o_0),
    .B2(n_6228_o_0),
    .Y(n_6382_o_0));
 OAI21xp33_ASAP7_75t_R n_6383 (.A1(n_6142_o_0),
    .A2(n_6382_o_0),
    .B(n_6075_o_0),
    .Y(n_6383_o_0));
 AO21x1_ASAP7_75t_R n_6384 (.A1(n_6128_o_0),
    .A2(n_6056_o_0),
    .B(n_6195_o_0),
    .Y(n_6384_o_0));
 OAI211xp5_ASAP7_75t_R n_6385 (.A1(n_6067_o_0),
    .A2(n_6241_o_0),
    .B(n_6197_o_0),
    .C(n_6195_o_0),
    .Y(n_6385_o_0));
 AOI31xp33_ASAP7_75t_R n_6386 (.A1(n_6002_o_0),
    .A2(n_6384_o_0),
    .A3(n_6385_o_0),
    .B(n_6183_o_0),
    .Y(n_6386_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6387 (.A1(n_6380_o_0),
    .A2(n_6185_o_0),
    .B(n_6383_o_0),
    .C(n_6386_o_0),
    .Y(n_6387_o_0));
 OAI22xp33_ASAP7_75t_R n_6388 (.A1(n_6313_o_0),
    .A2(n_6164_o_0),
    .B1(n_6219_o_0),
    .B2(n_6124_o_0),
    .Y(n_6388_o_0));
 NOR3xp33_ASAP7_75t_R n_6389 (.A(n_6124_o_0),
    .B(n_6219_o_0),
    .C(n_6067_o_0),
    .Y(n_6389_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6390 (.A1(n_6388_o_0),
    .A2(n_6067_o_0),
    .B(n_6389_o_0),
    .C(n_6195_o_0),
    .Y(n_6390_o_0));
 NOR2xp33_ASAP7_75t_R n_6391 (.A(n_6031_o_0),
    .B(n_6055_o_0),
    .Y(n_6391_o_0));
 OAI21xp33_ASAP7_75t_R n_6392 (.A1(n_6039_o_0),
    .A2(n_6391_o_0),
    .B(n_6142_o_0),
    .Y(n_6392_o_0));
 AOI31xp33_ASAP7_75t_R n_6393 (.A1(n_6241_o_0),
    .A2(n_6039_o_0),
    .A3(n_6092_o_0),
    .B(n_6392_o_0),
    .Y(n_6393_o_0));
 INVx1_ASAP7_75t_R n_6394 (.A(n_6393_o_0),
    .Y(n_6394_o_0));
 AOI21xp33_ASAP7_75t_R n_6395 (.A1(n_6204_o_0),
    .A2(n_6153_o_0),
    .B(n_6067_o_0),
    .Y(n_6395_o_0));
 AOI21xp33_ASAP7_75t_R n_6396 (.A1(n_6039_o_0),
    .A2(n_6071_o_0),
    .B(n_6067_o_0),
    .Y(n_6396_o_0));
 AOI21xp33_ASAP7_75t_R n_6397 (.A1(n_6057_o_0),
    .A2(n_6055_o_0),
    .B(n_6396_o_0),
    .Y(n_6397_o_0));
 OAI21xp33_ASAP7_75t_R n_6398 (.A1(n_6185_o_0),
    .A2(n_6397_o_0),
    .B(n_6003_o_0),
    .Y(n_6398_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6399 (.A1(n_6203_o_0),
    .A2(n_6395_o_0),
    .B(n_6142_o_0),
    .C(n_6398_o_0),
    .Y(n_6399_o_0));
 AOI31xp33_ASAP7_75t_R n_6400 (.A1(n_6159_o_0),
    .A2(n_6390_o_0),
    .A3(n_6394_o_0),
    .B(n_6399_o_0),
    .Y(n_6400_o_0));
 AOI21xp33_ASAP7_75t_R n_6401 (.A1(n_6183_o_0),
    .A2(n_6400_o_0),
    .B(n_6104_o_0),
    .Y(n_6401_o_0));
 AOI21xp33_ASAP7_75t_R n_6402 (.A1(n_6353_o_0),
    .A2(n_6194_o_0),
    .B(n_6003_o_0),
    .Y(n_6402_o_0));
 OAI211xp5_ASAP7_75t_R n_6403 (.A1(n_6114_o_0),
    .A2(n_6039_o_0),
    .B(n_6197_o_0),
    .C(n_6003_o_0),
    .Y(n_6403_o_0));
 OAI21xp33_ASAP7_75t_R n_6404 (.A1(n_6216_o_0),
    .A2(n_6403_o_0),
    .B(n_6186_o_0),
    .Y(n_6404_o_0));
 NAND2xp33_ASAP7_75t_R n_6405 (.A(n_6039_o_0),
    .B(n_6030_o_0),
    .Y(n_6405_o_0));
 AOI31xp33_ASAP7_75t_R n_6406 (.A1(n_6071_o_0),
    .A2(n_6058_o_0),
    .A3(n_6055_o_0),
    .B(n_6075_o_0),
    .Y(n_6406_o_0));
 OAI21xp33_ASAP7_75t_R n_6407 (.A1(n_6405_o_0),
    .A2(n_6050_o_0),
    .B(n_6406_o_0),
    .Y(n_6407_o_0));
 AOI211xp5_ASAP7_75t_R n_6408 (.A1(n_6030_o_0),
    .A2(n_6086_o_0),
    .B(n_6302_o_0),
    .C(n_6055_o_0),
    .Y(n_6408_o_0));
 NAND2xp33_ASAP7_75t_R n_6409 (.A(n_6030_o_0),
    .B(n_6086_o_0),
    .Y(n_6409_o_0));
 AOI21xp33_ASAP7_75t_R n_6410 (.A1(n_6256_o_0),
    .A2(n_6409_o_0),
    .B(n_6159_o_0),
    .Y(n_6410_o_0));
 OAI21xp33_ASAP7_75t_R n_6411 (.A1(n_6219_o_0),
    .A2(n_6366_o_0),
    .B(n_6410_o_0),
    .Y(n_6411_o_0));
 OAI211xp5_ASAP7_75t_R n_6412 (.A1(n_6407_o_0),
    .A2(n_6408_o_0),
    .B(n_6411_o_0),
    .C(n_6185_o_0),
    .Y(n_6412_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6413 (.A1(n_6111_o_0),
    .A2(n_6402_o_0),
    .B(n_6404_o_0),
    .C(n_6412_o_0),
    .Y(n_6413_o_0));
 NOR3xp33_ASAP7_75t_R n_6414 (.A(n_6072_o_0),
    .B(n_6092_o_0),
    .C(n_6214_o_0),
    .Y(n_6414_o_0));
 NOR4xp25_ASAP7_75t_R n_6415 (.A(n_6414_o_0),
    .B(n_6379_o_0),
    .C(n_6186_o_0),
    .D(n_6002_o_0),
    .Y(n_6415_o_0));
 INVx1_ASAP7_75t_R n_6416 (.A(n_6284_o_0),
    .Y(n_6416_o_0));
 NOR4xp25_ASAP7_75t_R n_6417 (.A(n_6416_o_0),
    .B(n_6205_o_0),
    .C(n_6186_o_0),
    .D(n_6075_o_0),
    .Y(n_6417_o_0));
 OAI21xp33_ASAP7_75t_R n_6418 (.A1(n_6206_o_0),
    .A2(n_6072_o_0),
    .B(n_6195_o_0),
    .Y(n_6418_o_0));
 AOI211xp5_ASAP7_75t_R n_6419 (.A1(n_6030_o_0),
    .A2(n_6039_o_0),
    .B(n_6143_o_0),
    .C(n_6092_o_0),
    .Y(n_6419_o_0));
 AOI21xp33_ASAP7_75t_R n_6420 (.A1(n_6058_o_0),
    .A2(n_6147_o_0),
    .B(n_6159_o_0),
    .Y(n_6420_o_0));
 OAI211xp5_ASAP7_75t_R n_6421 (.A1(n_6050_o_0),
    .A2(n_6109_o_0),
    .B(n_6420_o_0),
    .C(n_6195_o_0),
    .Y(n_6421_o_0));
 OAI31xp33_ASAP7_75t_R n_6422 (.A1(n_6075_o_0),
    .A2(n_6418_o_0),
    .A3(n_6419_o_0),
    .B(n_6421_o_0),
    .Y(n_6422_o_0));
 OAI31xp33_ASAP7_75t_R n_6423 (.A1(n_6415_o_0),
    .A2(n_6417_o_0),
    .A3(n_6422_o_0),
    .B(n_6107_o_0),
    .Y(n_6423_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6424 (.A1(n_6107_o_0),
    .A2(n_6413_o_0),
    .B(n_6423_o_0),
    .C(n_6105_o_0),
    .Y(n_6424_o_0));
 AOI21xp33_ASAP7_75t_R n_6425 (.A1(n_6387_o_0),
    .A2(n_6401_o_0),
    .B(n_6424_o_0),
    .Y(n_6425_o_0));
 AO21x1_ASAP7_75t_R n_6426 (.A1(n_6218_o_0),
    .A2(n_6191_o_0),
    .B(n_6269_o_0),
    .Y(n_6426_o_0));
 NAND2xp33_ASAP7_75t_R n_6427 (.A(n_6003_o_0),
    .B(n_6197_o_0),
    .Y(n_6427_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6428 (.A1(n_6039_o_0),
    .A2(n_6062_o_0),
    .B(n_6396_o_0),
    .C(n_6427_o_0),
    .Y(n_6428_o_0));
 AOI211xp5_ASAP7_75t_R n_6429 (.A1(n_6426_o_0),
    .A2(n_6159_o_0),
    .B(n_6428_o_0),
    .C(n_6195_o_0),
    .Y(n_6429_o_0));
 OAI21xp33_ASAP7_75t_R n_6430 (.A1(n_6017_o_0),
    .A2(n_6062_o_0),
    .B(n_6251_o_0),
    .Y(n_6430_o_0));
 OAI31xp33_ASAP7_75t_R n_6431 (.A1(n_6050_o_0),
    .A2(n_6109_o_0),
    .A3(n_6207_o_0),
    .B(n_6430_o_0),
    .Y(n_6431_o_0));
 OAI21xp33_ASAP7_75t_R n_6432 (.A1(n_6062_o_0),
    .A2(n_6092_o_0),
    .B(n_6159_o_0),
    .Y(n_6432_o_0));
 OAI21xp33_ASAP7_75t_R n_6433 (.A1(n_6432_o_0),
    .A2(n_6379_o_0),
    .B(n_6186_o_0),
    .Y(n_6433_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6434 (.A1(n_6431_o_0),
    .A2(n_6003_o_0),
    .B(n_6433_o_0),
    .C(n_6096_o_0),
    .Y(n_6434_o_0));
 AOI21xp33_ASAP7_75t_R n_6435 (.A1(n_6058_o_0),
    .A2(n_6224_o_0),
    .B(n_6089_o_0),
    .Y(n_6435_o_0));
 OAI311xp33_ASAP7_75t_R n_6436 (.A1(n_6062_o_0),
    .A2(n_6039_o_0),
    .A3(n_6031_o_0),
    .B1(n_6092_o_0),
    .C1(n_6110_o_0),
    .Y(n_6436_o_0));
 OAI31xp33_ASAP7_75t_R n_6437 (.A1(n_6031_o_0),
    .A2(n_6050_o_0),
    .A3(n_6302_o_0),
    .B(n_6436_o_0),
    .Y(n_6437_o_0));
 OAI321xp33_ASAP7_75t_R n_6438 (.A1(n_6003_o_0),
    .A2(n_6435_o_0),
    .A3(n_6168_o_0),
    .B1(n_6437_o_0),
    .B2(n_6159_o_0),
    .C(n_6195_o_0),
    .Y(n_6438_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6439 (.A1(n_6058_o_0),
    .A2(n_6031_o_0),
    .B(n_6336_o_0),
    .C(n_6092_o_0),
    .Y(n_6439_o_0));
 INVx1_ASAP7_75t_R n_6440 (.A(n_6208_o_0),
    .Y(n_6440_o_0));
 OAI211xp5_ASAP7_75t_R n_6441 (.A1(n_6440_o_0),
    .A2(n_6092_o_0),
    .B(n_6219_o_0),
    .C(n_6075_o_0),
    .Y(n_6441_o_0));
 OAI311xp33_ASAP7_75t_R n_6442 (.A1(n_6075_o_0),
    .A2(n_6439_o_0),
    .A3(n_6068_o_0),
    .B1(n_6185_o_0),
    .C1(n_6441_o_0),
    .Y(n_6442_o_0));
 NAND3xp33_ASAP7_75t_R n_6443 (.A(n_6438_o_0),
    .B(n_6442_o_0),
    .C(n_6183_o_0),
    .Y(n_6443_o_0));
 OAI21xp33_ASAP7_75t_R n_6444 (.A1(n_6429_o_0),
    .A2(n_6434_o_0),
    .B(n_6443_o_0),
    .Y(n_6444_o_0));
 AO22x1_ASAP7_75t_R n_6445 (.A1(n_6381_o_0),
    .A2(n_6092_o_0),
    .B1(n_6218_o_0),
    .B2(n_6084_o_0),
    .Y(n_6445_o_0));
 NAND3xp33_ASAP7_75t_R n_6446 (.A(n_6166_o_0),
    .B(n_6299_o_0),
    .C(n_6092_o_0),
    .Y(n_6446_o_0));
 OAI211xp5_ASAP7_75t_R n_6447 (.A1(n_6110_o_0),
    .A2(n_6092_o_0),
    .B(n_6446_o_0),
    .C(n_6185_o_0),
    .Y(n_6447_o_0));
 OAI21xp33_ASAP7_75t_R n_6448 (.A1(n_6185_o_0),
    .A2(n_6445_o_0),
    .B(n_6447_o_0),
    .Y(n_6448_o_0));
 NAND2xp33_ASAP7_75t_R n_6449 (.A(n_6031_o_0),
    .B(n_6067_o_0),
    .Y(n_6449_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6450 (.A1(n_6055_o_0),
    .A2(n_6254_o_0),
    .B(n_6449_o_0),
    .C(n_6237_o_0),
    .Y(n_6450_o_0));
 OAI31xp33_ASAP7_75t_R n_6451 (.A1(n_6086_o_0),
    .A2(n_6302_o_0),
    .A3(n_6055_o_0),
    .B(n_6142_o_0),
    .Y(n_6451_o_0));
 AO21x1_ASAP7_75t_R n_6452 (.A1(n_6165_o_0),
    .A2(n_6166_o_0),
    .B(n_6451_o_0),
    .Y(n_6452_o_0));
 OAI211xp5_ASAP7_75t_R n_6453 (.A1(n_6185_o_0),
    .A2(n_6450_o_0),
    .B(n_6452_o_0),
    .C(n_6159_o_0),
    .Y(n_6453_o_0));
 OAI21xp33_ASAP7_75t_R n_6454 (.A1(n_6002_o_0),
    .A2(n_6448_o_0),
    .B(n_6453_o_0),
    .Y(n_6454_o_0));
 INVx1_ASAP7_75t_R n_6455 (.A(n_6089_o_0),
    .Y(n_6455_o_0));
 OAI31xp33_ASAP7_75t_R n_6456 (.A1(n_6455_o_0),
    .A2(n_6216_o_0),
    .A3(n_6185_o_0),
    .B(n_6003_o_0),
    .Y(n_6456_o_0));
 OAI31xp33_ASAP7_75t_R n_6457 (.A1(n_6120_o_0),
    .A2(n_6088_o_0),
    .A3(n_6050_o_0),
    .B(n_6142_o_0),
    .Y(n_6457_o_0));
 AOI21xp33_ASAP7_75t_R n_6458 (.A1(n_6157_o_0),
    .A2(n_6299_o_0),
    .B(n_6457_o_0),
    .Y(n_6458_o_0));
 NAND3xp33_ASAP7_75t_R n_6459 (.A(n_6084_o_0),
    .B(n_6166_o_0),
    .C(n_6092_o_0),
    .Y(n_6459_o_0));
 INVx1_ASAP7_75t_R n_6460 (.A(n_6391_o_0),
    .Y(n_6460_o_0));
 AOI21xp33_ASAP7_75t_R n_6461 (.A1(n_6067_o_0),
    .A2(n_6114_o_0),
    .B(n_6195_o_0),
    .Y(n_6461_o_0));
 AOI33xp33_ASAP7_75t_R n_6462 (.A1(n_6186_o_0),
    .A2(n_6459_o_0),
    .A3(n_6324_o_0),
    .B1(n_6460_o_0),
    .B2(n_6461_o_0),
    .B3(n_6125_o_0),
    .Y(n_6462_o_0));
 AOI21xp33_ASAP7_75t_R n_6463 (.A1(n_6159_o_0),
    .A2(n_6462_o_0),
    .B(n_6107_o_0),
    .Y(n_6463_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6464 (.A1(n_6456_o_0),
    .A2(n_6458_o_0),
    .B(n_6463_o_0),
    .C(n_6104_o_0),
    .Y(n_6464_o_0));
 OAI21xp33_ASAP7_75t_R n_6465 (.A1(n_6096_o_0),
    .A2(n_6454_o_0),
    .B(n_6464_o_0),
    .Y(n_6465_o_0));
 OAI21xp33_ASAP7_75t_R n_6466 (.A1(n_6133_o_0),
    .A2(n_6444_o_0),
    .B(n_6465_o_0),
    .Y(n_6466_o_0));
 AO21x1_ASAP7_75t_R n_6467 (.A1(n_6191_o_0),
    .A2(n_6157_o_0),
    .B(n_6003_o_0),
    .Y(n_6467_o_0));
 AOI31xp33_ASAP7_75t_R n_6468 (.A1(n_6067_o_0),
    .A2(n_6084_o_0),
    .A3(n_6173_o_0),
    .B(n_6467_o_0),
    .Y(n_6468_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6469 (.A1(n_6067_o_0),
    .A2(n_6338_o_0),
    .B(n_6308_o_0),
    .C(n_6159_o_0),
    .Y(n_6469_o_0));
 AOI211xp5_ASAP7_75t_R n_6470 (.A1(n_6058_o_0),
    .A2(n_6031_o_0),
    .B(n_6124_o_0),
    .C(n_6055_o_0),
    .Y(n_6470_o_0));
 AOI211xp5_ASAP7_75t_R n_6471 (.A1(n_6030_o_0),
    .A2(n_6086_o_0),
    .B(n_6041_o_0),
    .C(n_6050_o_0),
    .Y(n_6471_o_0));
 OAI21xp33_ASAP7_75t_R n_6472 (.A1(n_6062_o_0),
    .A2(n_6254_o_0),
    .B(n_6055_o_0),
    .Y(n_6472_o_0));
 OAI211xp5_ASAP7_75t_R n_6473 (.A1(n_6110_o_0),
    .A2(n_6067_o_0),
    .B(n_6472_o_0),
    .C(n_6003_o_0),
    .Y(n_6473_o_0));
 OAI311xp33_ASAP7_75t_R n_6474 (.A1(n_6003_o_0),
    .A2(n_6470_o_0),
    .A3(n_6471_o_0),
    .B1(n_6142_o_0),
    .C1(n_6473_o_0),
    .Y(n_6474_o_0));
 OAI31xp33_ASAP7_75t_R n_6475 (.A1(n_6142_o_0),
    .A2(n_6468_o_0),
    .A3(n_6469_o_0),
    .B(n_6474_o_0),
    .Y(n_6475_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6476 (.A1(n_6031_o_0),
    .A2(n_6058_o_0),
    .B(n_6030_o_0),
    .C(n_6325_o_0),
    .Y(n_6476_o_0));
 INVx1_ASAP7_75t_R n_6477 (.A(n_6476_o_0),
    .Y(n_6477_o_0));
 OAI22xp33_ASAP7_75t_R n_6478 (.A1(n_6193_o_0),
    .A2(n_6109_o_0),
    .B1(n_6050_o_0),
    .B2(n_6477_o_0),
    .Y(n_6478_o_0));
 OAI31xp33_ASAP7_75t_R n_6479 (.A1(n_6058_o_0),
    .A2(n_6065_o_0),
    .A3(n_6067_o_0),
    .B(n_6003_o_0),
    .Y(n_6479_o_0));
 AOI21xp33_ASAP7_75t_R n_6480 (.A1(n_6017_o_0),
    .A2(n_6039_o_0),
    .B(n_6267_o_0),
    .Y(n_6480_o_0));
 AOI211xp5_ASAP7_75t_R n_6481 (.A1(n_6050_o_0),
    .A2(n_6254_o_0),
    .B(n_6479_o_0),
    .C(n_6480_o_0),
    .Y(n_6481_o_0));
 AOI21xp33_ASAP7_75t_R n_6482 (.A1(n_6159_o_0),
    .A2(n_6478_o_0),
    .B(n_6481_o_0),
    .Y(n_6482_o_0));
 OAI321xp33_ASAP7_75t_R n_6483 (.A1(n_6092_o_0),
    .A2(n_6227_o_0),
    .A3(n_6202_o_0),
    .B1(n_6030_o_0),
    .B2(n_6067_o_0),
    .C(n_6159_o_0),
    .Y(n_6483_o_0));
 NAND4xp25_ASAP7_75t_R n_6484 (.A(n_6055_o_0),
    .B(n_6062_o_0),
    .C(n_6017_o_0),
    .D(n_6039_o_0),
    .Y(n_6484_o_0));
 NAND4xp25_ASAP7_75t_R n_6485 (.A(n_6336_o_0),
    .B(n_6484_o_0),
    .C(n_6315_o_0),
    .D(n_6003_o_0),
    .Y(n_6485_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6486 (.A1(n_6483_o_0),
    .A2(n_6485_o_0),
    .B(n_6142_o_0),
    .C(n_6107_o_0),
    .Y(n_6486_o_0));
 AOI21xp33_ASAP7_75t_R n_6487 (.A1(n_6142_o_0),
    .A2(n_6482_o_0),
    .B(n_6486_o_0),
    .Y(n_6487_o_0));
 AOI21xp33_ASAP7_75t_R n_6488 (.A1(n_6096_o_0),
    .A2(n_6475_o_0),
    .B(n_6487_o_0),
    .Y(n_6488_o_0));
 OAI31xp33_ASAP7_75t_R n_6489 (.A1(n_6086_o_0),
    .A2(n_6085_o_0),
    .A3(n_6055_o_0),
    .B(n_6075_o_0),
    .Y(n_6489_o_0));
 AOI21xp33_ASAP7_75t_R n_6490 (.A1(n_6067_o_0),
    .A2(n_6156_o_0),
    .B(n_6489_o_0),
    .Y(n_6490_o_0));
 INVx1_ASAP7_75t_R n_6491 (.A(n_6157_o_0),
    .Y(n_6491_o_0));
 OAI21xp33_ASAP7_75t_R n_6492 (.A1(n_6114_o_0),
    .A2(n_6039_o_0),
    .B(n_6165_o_0),
    .Y(n_6492_o_0));
 AOI21xp33_ASAP7_75t_R n_6493 (.A1(n_6491_o_0),
    .A2(n_6492_o_0),
    .B(n_6075_o_0),
    .Y(n_6493_o_0));
 OAI21xp33_ASAP7_75t_R n_6494 (.A1(n_6050_o_0),
    .A2(n_6237_o_0),
    .B(n_6193_o_0),
    .Y(n_6494_o_0));
 NAND2xp33_ASAP7_75t_R n_6495 (.A(n_6062_o_0),
    .B(n_6449_o_0),
    .Y(n_6495_o_0));
 AOI31xp33_ASAP7_75t_R n_6496 (.A1(n_6053_o_0),
    .A2(n_6495_o_0),
    .A3(n_6002_o_0),
    .B(n_6142_o_0),
    .Y(n_6496_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6497 (.A1(n_6040_o_0),
    .A2(n_6494_o_0),
    .B(n_6159_o_0),
    .C(n_6496_o_0),
    .Y(n_6497_o_0));
 OAI31xp33_ASAP7_75t_R n_6498 (.A1(n_6186_o_0),
    .A2(n_6490_o_0),
    .A3(n_6493_o_0),
    .B(n_6497_o_0),
    .Y(n_6498_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6499 (.A1(n_6215_o_0),
    .A2(n_6405_o_0),
    .B(n_6050_o_0),
    .C(n_6002_o_0),
    .Y(n_6499_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6500 (.A1(n_6065_o_0),
    .A2(n_6039_o_0),
    .B(n_6455_o_0),
    .C(n_6159_o_0),
    .Y(n_6500_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6501 (.A1(n_6053_o_0),
    .A2(n_6055_o_0),
    .B(n_6500_o_0),
    .C(n_6142_o_0),
    .Y(n_6501_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6502 (.A1(n_6381_o_0),
    .A2(n_6092_o_0),
    .B(n_6499_o_0),
    .C(n_6501_o_0),
    .Y(n_6502_o_0));
 OAI211xp5_ASAP7_75t_R n_6503 (.A1(n_6030_o_0),
    .A2(n_6039_o_0),
    .B(n_6110_o_0),
    .C(n_6067_o_0),
    .Y(n_6503_o_0));
 AOI31xp33_ASAP7_75t_R n_6504 (.A1(n_6075_o_0),
    .A2(n_6503_o_0),
    .A3(n_6115_o_0),
    .B(n_6186_o_0),
    .Y(n_6504_o_0));
 OAI21xp33_ASAP7_75t_R n_6505 (.A1(n_6003_o_0),
    .A2(n_6303_o_0),
    .B(n_6504_o_0),
    .Y(n_6505_o_0));
 AOI31xp33_ASAP7_75t_R n_6506 (.A1(n_5995_o_0),
    .A2(n_6502_o_0),
    .A3(n_6505_o_0),
    .B(n_6104_o_0),
    .Y(n_6506_o_0));
 OAI21xp33_ASAP7_75t_R n_6507 (.A1(n_6096_o_0),
    .A2(n_6498_o_0),
    .B(n_6506_o_0),
    .Y(n_6507_o_0));
 OAI21xp33_ASAP7_75t_R n_6508 (.A1(n_6133_o_0),
    .A2(n_6488_o_0),
    .B(n_6507_o_0),
    .Y(n_6508_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6509 (.A1(n_6039_o_0),
    .A2(n_6017_o_0),
    .B(n_6030_o_0),
    .C(n_6067_o_0),
    .Y(n_6509_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6510 (.A1(n_6031_o_0),
    .A2(n_6030_o_0),
    .B(n_6050_o_0),
    .C(n_6148_o_0),
    .Y(n_6510_o_0));
 OAI31xp33_ASAP7_75t_R n_6511 (.A1(n_6002_o_0),
    .A2(n_6203_o_0),
    .A3(n_6509_o_0),
    .B(n_6510_o_0),
    .Y(n_6511_o_0));
 NOR2xp33_ASAP7_75t_R n_6512 (.A(n_6039_o_0),
    .B(n_6065_o_0),
    .Y(n_6512_o_0));
 OAI22xp33_ASAP7_75t_R n_6513 (.A1(n_6512_o_0),
    .A2(n_6242_o_0),
    .B1(n_6082_o_0),
    .B2(n_6214_o_0),
    .Y(n_6513_o_0));
 OAI21xp33_ASAP7_75t_R n_6514 (.A1(n_6030_o_0),
    .A2(n_6058_o_0),
    .B(n_6067_o_0),
    .Y(n_6514_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6515 (.A1(n_6065_o_0),
    .A2(n_6039_o_0),
    .B(n_6055_o_0),
    .C(n_6514_o_0),
    .Y(n_6515_o_0));
 INVx1_ASAP7_75t_R n_6516 (.A(n_6179_o_0),
    .Y(n_6516_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6517 (.A1(n_6515_o_0),
    .A2(n_6516_o_0),
    .B(n_6003_o_0),
    .C(n_6185_o_0),
    .Y(n_6517_o_0));
 AOI21xp33_ASAP7_75t_R n_6518 (.A1(n_6075_o_0),
    .A2(n_6513_o_0),
    .B(n_6517_o_0),
    .Y(n_6518_o_0));
 AOI21xp33_ASAP7_75t_R n_6519 (.A1(n_6195_o_0),
    .A2(n_6511_o_0),
    .B(n_6518_o_0),
    .Y(n_6519_o_0));
 INVx1_ASAP7_75t_R n_6520 (.A(n_6251_o_0),
    .Y(n_6520_o_0));
 NAND2xp33_ASAP7_75t_R n_6521 (.A(n_6110_o_0),
    .B(n_6218_o_0),
    .Y(n_6521_o_0));
 OAI31xp33_ASAP7_75t_R n_6522 (.A1(n_6223_o_0),
    .A2(n_6266_o_0),
    .A3(n_6520_o_0),
    .B(n_6521_o_0),
    .Y(n_6522_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6523 (.A1(n_6017_o_0),
    .A2(n_6062_o_0),
    .B(n_6239_o_0),
    .C(n_6159_o_0),
    .Y(n_6523_o_0));
 AO21x1_ASAP7_75t_R n_6524 (.A1(n_6523_o_0),
    .A2(n_6332_o_0),
    .B(n_6185_o_0),
    .Y(n_6524_o_0));
 OAI221xp5_ASAP7_75t_R n_6525 (.A1(n_6092_o_0),
    .A2(n_6204_o_0),
    .B1(n_6147_o_0),
    .B2(n_6039_o_0),
    .C(n_6148_o_0),
    .Y(n_6525_o_0));
 AOI31xp33_ASAP7_75t_R n_6526 (.A1(n_6052_o_0),
    .A2(n_6278_o_0),
    .A3(n_6055_o_0),
    .B(n_6002_o_0),
    .Y(n_6526_o_0));
 OAI21xp33_ASAP7_75t_R n_6527 (.A1(n_6067_o_0),
    .A2(n_6224_o_0),
    .B(n_6526_o_0),
    .Y(n_6527_o_0));
 NAND3xp33_ASAP7_75t_R n_6528 (.A(n_6525_o_0),
    .B(n_6527_o_0),
    .C(n_6142_o_0),
    .Y(n_6528_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6529 (.A1(n_6522_o_0),
    .A2(n_6159_o_0),
    .B(n_6524_o_0),
    .C(n_6528_o_0),
    .Y(n_6529_o_0));
 OAI22xp33_ASAP7_75t_R n_6530 (.A1(n_6519_o_0),
    .A2(n_6183_o_0),
    .B1(n_6529_o_0),
    .B2(n_5995_o_0),
    .Y(n_6530_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6531 (.A1(n_6325_o_0),
    .A2(n_6068_o_0),
    .B(n_6243_o_0),
    .C(n_6142_o_0),
    .Y(n_6531_o_0));
 AOI21xp33_ASAP7_75t_R n_6532 (.A1(n_6204_o_0),
    .A2(n_6153_o_0),
    .B(n_6092_o_0),
    .Y(n_6532_o_0));
 AOI21xp33_ASAP7_75t_R n_6533 (.A1(n_6173_o_0),
    .A2(n_6391_o_0),
    .B(n_6165_o_0),
    .Y(n_6533_o_0));
 OAI21xp33_ASAP7_75t_R n_6534 (.A1(n_6532_o_0),
    .A2(n_6533_o_0),
    .B(n_6186_o_0),
    .Y(n_6534_o_0));
 AOI31xp33_ASAP7_75t_R n_6535 (.A1(n_6192_o_0),
    .A2(n_6110_o_0),
    .A3(n_6092_o_0),
    .B(n_6075_o_0),
    .Y(n_6535_o_0));
 OAI21xp33_ASAP7_75t_R n_6536 (.A1(n_6195_o_0),
    .A2(n_6279_o_0),
    .B(n_6535_o_0),
    .Y(n_6536_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6537 (.A1(n_6381_o_0),
    .A2(n_6067_o_0),
    .B(n_6194_o_0),
    .C(n_6195_o_0),
    .D(n_6536_o_0),
    .Y(n_6537_o_0));
 AOI31xp33_ASAP7_75t_R n_6538 (.A1(n_6003_o_0),
    .A2(n_6531_o_0),
    .A3(n_6534_o_0),
    .B(n_6537_o_0),
    .Y(n_6538_o_0));
 OAI21xp33_ASAP7_75t_R n_6539 (.A1(n_5995_o_0),
    .A2(n_6538_o_0),
    .B(n_6133_o_0),
    .Y(n_6539_o_0));
 NOR2xp33_ASAP7_75t_R n_6540 (.A(n_6050_o_0),
    .B(n_6207_o_0),
    .Y(n_6540_o_0));
 INVx1_ASAP7_75t_R n_6541 (.A(n_6293_o_0),
    .Y(n_6541_o_0));
 NAND2xp33_ASAP7_75t_R n_6542 (.A(n_6108_o_0),
    .B(n_6238_o_0),
    .Y(n_6542_o_0));
 OAI31xp33_ASAP7_75t_R n_6543 (.A1(n_6055_o_0),
    .A2(n_6541_o_0),
    .A3(n_6172_o_0),
    .B(n_6542_o_0),
    .Y(n_6543_o_0));
 AOI21xp33_ASAP7_75t_R n_6544 (.A1(n_6195_o_0),
    .A2(n_6543_o_0),
    .B(n_6003_o_0),
    .Y(n_6544_o_0));
 OAI31xp33_ASAP7_75t_R n_6545 (.A1(n_6068_o_0),
    .A2(n_6186_o_0),
    .A3(n_6540_o_0),
    .B(n_6544_o_0),
    .Y(n_6545_o_0));
 OAI211xp5_ASAP7_75t_R n_6546 (.A1(n_6065_o_0),
    .A2(n_6039_o_0),
    .B(n_6092_o_0),
    .C(n_6293_o_0),
    .Y(n_6546_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6547 (.A1(n_6030_o_0),
    .A2(n_6086_o_0),
    .B(n_6050_o_0),
    .C(n_6546_o_0),
    .Y(n_6547_o_0));
 AOI21xp33_ASAP7_75t_R n_6548 (.A1(n_6185_o_0),
    .A2(n_6547_o_0),
    .B(n_6159_o_0),
    .Y(n_6548_o_0));
 OAI31xp33_ASAP7_75t_R n_6549 (.A1(n_6185_o_0),
    .A2(n_6391_o_0),
    .A3(n_6419_o_0),
    .B(n_6548_o_0),
    .Y(n_6549_o_0));
 AOI21xp33_ASAP7_75t_R n_6550 (.A1(n_6545_o_0),
    .A2(n_6549_o_0),
    .B(n_6107_o_0),
    .Y(n_6550_o_0));
 OAI22xp33_ASAP7_75t_R n_6551 (.A1(n_6530_o_0),
    .A2(n_6105_o_0),
    .B1(n_6539_o_0),
    .B2(n_6550_o_0),
    .Y(n_6551_o_0));
 XNOR2xp5_ASAP7_75t_R n_6552 (.A(_01017_),
    .B(_01056_),
    .Y(n_6552_o_0));
 XNOR2xp5_ASAP7_75t_R n_6553 (.A(_01064_),
    .B(n_6552_o_0),
    .Y(n_6553_o_0));
 XOR2xp5_ASAP7_75t_R n_6554 (.A(n_4298_o_0),
    .B(n_6553_o_0),
    .Y(n_6554_o_0));
 NOR2xp33_ASAP7_75t_R n_6555 (.A(_00696_),
    .B(net),
    .Y(n_6555_o_0));
 AOI21xp33_ASAP7_75t_R n_6556 (.A1(net),
    .A2(n_6554_o_0),
    .B(n_6555_o_0),
    .Y(n_6556_o_0));
 XOR2xp5_ASAP7_75t_R n_6557 (.A(_00945_),
    .B(n_6556_o_0),
    .Y(n_6557_o_0));
 INVx1_ASAP7_75t_R n_6558 (.A(n_6557_o_0),
    .Y(n_6558_o_0));
 XNOR2xp5_ASAP7_75t_R n_6559 (.A(_01066_),
    .B(_01067_),
    .Y(n_6559_o_0));
 XNOR2xp5_ASAP7_75t_R n_6560 (.A(_01106_),
    .B(n_6559_o_0),
    .Y(n_6560_o_0));
 XOR2xp5_ASAP7_75t_R n_6561 (.A(_01019_),
    .B(_01058_),
    .Y(n_6561_o_0));
 NOR2xp33_ASAP7_75t_R n_6562 (.A(n_6561_o_0),
    .B(n_6560_o_0),
    .Y(n_6562_o_0));
 NOR2xp33_ASAP7_75t_R n_6563 (.A(_00694_),
    .B(net),
    .Y(n_6563_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6564 (.A1(n_6560_o_0),
    .A2(n_6561_o_0),
    .B(n_6562_o_0),
    .C(net),
    .D(n_6563_o_0),
    .Y(n_6564_o_0));
 XNOR2xp5_ASAP7_75t_R n_6565 (.A(_00947_),
    .B(n_6564_o_0),
    .Y(n_6565_o_0));
 INVx1_ASAP7_75t_R n_6566 (.A(n_6565_o_0),
    .Y(n_6566_o_0));
 XNOR2xp5_ASAP7_75t_R n_6567 (.A(_01016_),
    .B(n_4265_o_0),
    .Y(n_6567_o_0));
 XNOR2xp5_ASAP7_75t_R n_6568 (.A(_01063_),
    .B(_01067_),
    .Y(n_6568_o_0));
 XNOR2xp5_ASAP7_75t_R n_6569 (.A(n_4266_o_0),
    .B(n_6568_o_0),
    .Y(n_6569_o_0));
 XNOR2xp5_ASAP7_75t_R n_6570 (.A(n_6567_o_0),
    .B(n_6569_o_0),
    .Y(n_6570_o_0));
 OR2x2_ASAP7_75t_R n_6571 (.A(_00697_),
    .B(net),
    .Y(n_6571_o_0));
 OAI21xp33_ASAP7_75t_R n_6572 (.A1(net9),
    .A2(n_6570_o_0),
    .B(n_6571_o_0),
    .Y(n_6572_o_0));
 XNOR2xp5_ASAP7_75t_R n_6573 (.A(_00944_),
    .B(n_6572_o_0),
    .Y(n_6573_o_0));
 XNOR2xp5_ASAP7_75t_R n_6574 (.A(_01060_),
    .B(_01067_),
    .Y(n_6574_o_0));
 INVx1_ASAP7_75t_R n_6575 (.A(n_6574_o_0),
    .Y(n_6575_o_0));
 XOR2xp5_ASAP7_75t_R n_6576 (.A(_01059_),
    .B(_01099_),
    .Y(n_6576_o_0));
 INVx1_ASAP7_75t_R n_6577 (.A(_01012_),
    .Y(n_6577_o_0));
 NAND2xp33_ASAP7_75t_R n_6578 (.A(n_6577_o_0),
    .B(n_6576_o_0),
    .Y(n_6578_o_0));
 OAI21xp33_ASAP7_75t_R n_6579 (.A1(n_6576_o_0),
    .A2(n_6577_o_0),
    .B(n_6578_o_0),
    .Y(n_6579_o_0));
 NOR2xp33_ASAP7_75t_R n_6580 (.A(n_6577_o_0),
    .B(n_6576_o_0),
    .Y(n_6580_o_0));
 AOI211xp5_ASAP7_75t_R n_6581 (.A1(n_6576_o_0),
    .A2(n_6577_o_0),
    .B(n_6580_o_0),
    .C(n_6575_o_0),
    .Y(n_6581_o_0));
 NOR2xp33_ASAP7_75t_R n_6582 (.A(_00550_),
    .B(_00858_),
    .Y(n_6582_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6583 (.A1(n_6575_o_0),
    .A2(n_6579_o_0),
    .B(n_6581_o_0),
    .C(net77),
    .D(n_6582_o_0),
    .Y(n_6583_o_0));
 OAI211xp5_ASAP7_75t_R n_6584 (.A1(n_6576_o_0),
    .A2(n_6577_o_0),
    .B(n_6578_o_0),
    .C(n_6574_o_0),
    .Y(n_6584_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6585 (.A1(n_6576_o_0),
    .A2(n_6577_o_0),
    .B(n_6580_o_0),
    .C(n_6575_o_0),
    .Y(n_6585_o_0));
 INVx1_ASAP7_75t_R n_6586 (.A(n_6582_o_0),
    .Y(n_6586_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6587 (.A1(n_6584_o_0),
    .A2(n_6585_o_0),
    .B(net1),
    .C(n_6586_o_0),
    .D(_00940_),
    .Y(n_6587_o_0));
 AO21x1_ASAP7_75t_R n_6588 (.A1(_00940_),
    .A2(n_6583_o_0),
    .B(n_6587_o_0),
    .Y(n_6588_o_0));
 XOR2xp5_ASAP7_75t_R n_6589 (.A(_01061_),
    .B(_01100_),
    .Y(n_6589_o_0));
 XNOR2xp5_ASAP7_75t_R n_6590 (.A(n_6574_o_0),
    .B(n_6589_o_0),
    .Y(n_6590_o_0));
 XNOR2xp5_ASAP7_75t_R n_6591 (.A(_01013_),
    .B(n_4205_o_0),
    .Y(n_6591_o_0));
 NOR2xp33_ASAP7_75t_R n_6592 (.A(n_6591_o_0),
    .B(n_6590_o_0),
    .Y(n_6592_o_0));
 NOR2xp33_ASAP7_75t_R n_6593 (.A(_00549_),
    .B(_00858_),
    .Y(n_6593_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6594 (.A1(n_6590_o_0),
    .A2(n_6591_o_0),
    .B(n_6592_o_0),
    .C(net77),
    .D(n_6593_o_0),
    .Y(n_6594_o_0));
 NOR2xp33_ASAP7_75t_R n_6595 (.A(_01013_),
    .B(n_4209_o_0),
    .Y(n_6595_o_0));
 XOR2xp5_ASAP7_75t_R n_6596 (.A(n_6574_o_0),
    .B(n_6589_o_0),
    .Y(n_6596_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6597 (.A1(_01013_),
    .A2(n_4209_o_0),
    .B(n_6595_o_0),
    .C(n_6596_o_0),
    .Y(n_6597_o_0));
 NAND2xp33_ASAP7_75t_R n_6598 (.A(n_6591_o_0),
    .B(n_6590_o_0),
    .Y(n_6598_o_0));
 INVx1_ASAP7_75t_R n_6599 (.A(n_6593_o_0),
    .Y(n_6599_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6600 (.A1(n_6597_o_0),
    .A2(n_6598_o_0),
    .B(net5),
    .C(n_6599_o_0),
    .D(_00941_),
    .Y(n_6600_o_0));
 AOI21xp5_ASAP7_75t_R n_6601 (.A1(_00941_),
    .A2(n_6594_o_0),
    .B(n_6600_o_0),
    .Y(n_6601_o_0));
 NAND2xp33_ASAP7_75t_R n_6602 (.A(n_6588_o_0),
    .B(n_6601_o_0),
    .Y(n_6602_o_0));
 AOI21x1_ASAP7_75t_R n_6603 (.A1(_00940_),
    .A2(n_6583_o_0),
    .B(n_6587_o_0),
    .Y(n_6603_o_0));
 INVx1_ASAP7_75t_R n_6604 (.A(_00942_),
    .Y(n_6604_o_0));
 NAND2xp33_ASAP7_75t_R n_6605 (.A(_01014_),
    .B(n_4186_o_0),
    .Y(n_6605_o_0));
 OAI21xp33_ASAP7_75t_R n_6606 (.A1(_01014_),
    .A2(n_4186_o_0),
    .B(n_6605_o_0),
    .Y(n_6606_o_0));
 OAI211xp5_ASAP7_75t_R n_6607 (.A1(_01014_),
    .A2(n_4186_o_0),
    .B(n_6605_o_0),
    .C(n_4210_o_0),
    .Y(n_6607_o_0));
 INVx1_ASAP7_75t_R n_6608 (.A(n_6607_o_0),
    .Y(n_6608_o_0));
 NOR2xp33_ASAP7_75t_R n_6609 (.A(_00552_),
    .B(net39),
    .Y(n_6609_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6610 (.A1(n_4206_o_0),
    .A2(n_6606_o_0),
    .B(n_6608_o_0),
    .C(net39),
    .D(n_6609_o_0),
    .Y(n_6610_o_0));
 NAND2xp33_ASAP7_75t_R n_6611 (.A(n_4206_o_0),
    .B(n_6606_o_0),
    .Y(n_6611_o_0));
 INVx1_ASAP7_75t_R n_6612 (.A(n_6609_o_0),
    .Y(n_6612_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6613 (.A1(n_6607_o_0),
    .A2(n_6611_o_0),
    .B(n_3021_o_0),
    .C(n_6612_o_0),
    .D(n_6604_o_0),
    .Y(n_6613_o_0));
 AOI21x1_ASAP7_75t_R n_6614 (.A1(n_6604_o_0),
    .A2(n_6610_o_0),
    .B(n_6613_o_0),
    .Y(n_6614_o_0));
 NAND2xp33_ASAP7_75t_R n_6615 (.A(n_6603_o_0),
    .B(n_6614_o_0),
    .Y(n_6615_o_0));
 XNOR2xp5_ASAP7_75t_R n_6616 (.A(_01062_),
    .B(_01067_),
    .Y(n_6616_o_0));
 XNOR2xp5_ASAP7_75t_R n_6617 (.A(n_4249_o_0),
    .B(n_6616_o_0),
    .Y(n_6617_o_0));
 XOR2xp5_ASAP7_75t_R n_6618 (.A(_01015_),
    .B(n_4248_o_0),
    .Y(n_6618_o_0));
 NAND2xp33_ASAP7_75t_R n_6619 (.A(n_6617_o_0),
    .B(n_6618_o_0),
    .Y(n_6619_o_0));
 OAI21xp33_ASAP7_75t_R n_6620 (.A1(n_6617_o_0),
    .A2(n_6618_o_0),
    .B(n_6619_o_0),
    .Y(n_6620_o_0));
 NOR2xp33_ASAP7_75t_R n_6621 (.A(_00698_),
    .B(_00858_),
    .Y(n_6621_o_0));
 AO21x1_ASAP7_75t_R n_6622 (.A1(n_6620_o_0),
    .A2(net39),
    .B(n_6621_o_0),
    .Y(n_6622_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6623 (.A1(n_6620_o_0),
    .A2(net),
    .B(n_6621_o_0),
    .C(_00943_),
    .Y(n_6623_o_0));
 OAI21x1_ASAP7_75t_R n_6624 (.A1(_00943_),
    .A2(n_6622_o_0),
    .B(n_6623_o_0),
    .Y(n_6624_o_0));
 NAND3xp33_ASAP7_75t_R n_6625 (.A(n_6602_o_0),
    .B(n_6615_o_0),
    .C(n_6624_o_0),
    .Y(n_6625_o_0));
 NAND2xp33_ASAP7_75t_R n_6626 (.A(n_6573_o_0),
    .B(n_6625_o_0),
    .Y(n_6626_o_0));
 INVx1_ASAP7_75t_R n_6627 (.A(n_6626_o_0),
    .Y(n_6627_o_0));
 AO21x1_ASAP7_75t_R n_6628 (.A1(n_6594_o_0),
    .A2(_00941_),
    .B(n_6600_o_0),
    .Y(n_6628_o_0));
 NAND2xp33_ASAP7_75t_R n_6629 (.A(n_6588_o_0),
    .B(n_6628_o_0),
    .Y(n_6629_o_0));
 AO21x2_ASAP7_75t_R n_6630 (.A1(n_6604_o_0),
    .A2(n_6610_o_0),
    .B(n_6613_o_0),
    .Y(n_6630_o_0));
 INVx1_ASAP7_75t_R n_6631 (.A(_00943_),
    .Y(n_6631_o_0));
 AOI211xp5_ASAP7_75t_R n_6632 (.A1(n_6620_o_0),
    .A2(net),
    .B(n_6631_o_0),
    .C(n_6621_o_0),
    .Y(n_6632_o_0));
 AOI21xp33_ASAP7_75t_R n_6633 (.A1(n_6631_o_0),
    .A2(n_6622_o_0),
    .B(n_6632_o_0),
    .Y(n_6633_o_0));
 AOI21xp33_ASAP7_75t_R n_6634 (.A1(n_6630_o_0),
    .A2(n_6603_o_0),
    .B(n_6633_o_0),
    .Y(n_6634_o_0));
 NAND2xp33_ASAP7_75t_R n_6635 (.A(n_6629_o_0),
    .B(n_6634_o_0),
    .Y(n_6635_o_0));
 NOR2xp33_ASAP7_75t_R n_6636 (.A(n_6628_o_0),
    .B(n_6615_o_0),
    .Y(n_6636_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6637 (.A1(_00941_),
    .A2(n_6594_o_0),
    .B(n_6600_o_0),
    .C(n_6588_o_0),
    .Y(n_6637_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6638 (.A1(n_6590_o_0),
    .A2(n_6591_o_0),
    .B(n_6592_o_0),
    .C(net),
    .Y(n_6638_o_0));
 OAI211xp5_ASAP7_75t_R n_6639 (.A1(_00549_),
    .A2(net),
    .B(n_6638_o_0),
    .C(_00941_),
    .Y(n_6639_o_0));
 OAI211xp5_ASAP7_75t_R n_6640 (.A1(_00941_),
    .A2(n_6594_o_0),
    .B(n_6639_o_0),
    .C(n_6603_o_0),
    .Y(n_6640_o_0));
 AOI21xp33_ASAP7_75t_R n_6641 (.A1(n_6637_o_0),
    .A2(n_6640_o_0),
    .B(n_6614_o_0),
    .Y(n_6641_o_0));
 NOR3xp33_ASAP7_75t_R n_6642 (.A(n_6636_o_0),
    .B(n_6641_o_0),
    .C(n_6633_o_0),
    .Y(n_6642_o_0));
 INVx1_ASAP7_75t_R n_6643 (.A(n_6600_o_0),
    .Y(n_6643_o_0));
 AOI21xp33_ASAP7_75t_R n_6644 (.A1(n_6643_o_0),
    .A2(n_6639_o_0),
    .B(n_6603_o_0),
    .Y(n_6644_o_0));
 NAND2xp33_ASAP7_75t_R n_6645 (.A(n_6614_o_0),
    .B(n_6644_o_0),
    .Y(n_6645_o_0));
 NAND3xp33_ASAP7_75t_R n_6646 (.A(n_6628_o_0),
    .B(n_6630_o_0),
    .C(n_6603_o_0),
    .Y(n_6646_o_0));
 AND3x1_ASAP7_75t_R n_6647 (.A(n_6645_o_0),
    .B(n_6646_o_0),
    .C(n_6624_o_0),
    .Y(n_6647_o_0));
 NAND2xp33_ASAP7_75t_R n_6648 (.A(_00944_),
    .B(n_6572_o_0),
    .Y(n_6648_o_0));
 OAI21xp5_ASAP7_75t_R n_6649 (.A1(_00944_),
    .A2(n_6572_o_0),
    .B(n_6648_o_0),
    .Y(n_6649_o_0));
 XNOR2xp5_ASAP7_75t_R n_6650 (.A(_01065_),
    .B(_01066_),
    .Y(n_6650_o_0));
 XNOR2xp5_ASAP7_75t_R n_6651 (.A(_01105_),
    .B(n_6650_o_0),
    .Y(n_6651_o_0));
 XOR2xp5_ASAP7_75t_R n_6652 (.A(_01018_),
    .B(_01057_),
    .Y(n_6652_o_0));
 NOR2xp33_ASAP7_75t_R n_6653 (.A(n_6652_o_0),
    .B(n_6651_o_0),
    .Y(n_6653_o_0));
 NOR2xp33_ASAP7_75t_R n_6654 (.A(_00695_),
    .B(net),
    .Y(n_6654_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6655 (.A1(n_6651_o_0),
    .A2(n_6652_o_0),
    .B(n_6653_o_0),
    .C(net),
    .D(n_6654_o_0),
    .Y(n_6655_o_0));
 NAND2xp33_ASAP7_75t_R n_6656 (.A(_00946_),
    .B(n_6655_o_0),
    .Y(n_6656_o_0));
 OAI21xp33_ASAP7_75t_R n_6657 (.A1(_00946_),
    .A2(n_6655_o_0),
    .B(n_6656_o_0),
    .Y(n_6657_o_0));
 OAI31xp33_ASAP7_75t_R n_6658 (.A1(n_6642_o_0),
    .A2(n_6647_o_0),
    .A3(n_6649_o_0),
    .B(n_6657_o_0),
    .Y(n_6658_o_0));
 XOR2xp5_ASAP7_75t_R n_6659 (.A(_00944_),
    .B(n_6572_o_0),
    .Y(n_6659_o_0));
 AOI211xp5_ASAP7_75t_R n_6660 (.A1(n_6620_o_0),
    .A2(net),
    .B(_00943_),
    .C(n_6621_o_0),
    .Y(n_6660_o_0));
 AOI21xp33_ASAP7_75t_R n_6661 (.A1(_00943_),
    .A2(n_6622_o_0),
    .B(n_6660_o_0),
    .Y(n_6661_o_0));
 AOI21xp33_ASAP7_75t_R n_6662 (.A1(n_6601_o_0),
    .A2(n_6603_o_0),
    .B(n_6630_o_0),
    .Y(n_6662_o_0));
 NAND3xp33_ASAP7_75t_R n_6663 (.A(n_6601_o_0),
    .B(n_6614_o_0),
    .C(n_6588_o_0),
    .Y(n_6663_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6664 (.A1(n_6610_o_0),
    .A2(n_6604_o_0),
    .B(n_6613_o_0),
    .C(n_6588_o_0),
    .Y(n_6664_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6665 (.A1(n_6620_o_0),
    .A2(net),
    .B(n_6621_o_0),
    .C(n_6631_o_0),
    .Y(n_6665_o_0));
 OAI21x1_ASAP7_75t_R n_6666 (.A1(n_6631_o_0),
    .A2(n_6622_o_0),
    .B(n_6665_o_0),
    .Y(n_6666_o_0));
 NAND3xp33_ASAP7_75t_R n_6667 (.A(n_6663_o_0),
    .B(n_6664_o_0),
    .C(n_6666_o_0),
    .Y(n_6667_o_0));
 OAI31xp33_ASAP7_75t_R n_6668 (.A1(n_6661_o_0),
    .A2(n_6641_o_0),
    .A3(n_6662_o_0),
    .B(n_6667_o_0),
    .Y(n_6668_o_0));
 INVx1_ASAP7_75t_R n_6669 (.A(n_6663_o_0),
    .Y(n_6669_o_0));
 OAI21xp33_ASAP7_75t_R n_6670 (.A1(n_6603_o_0),
    .A2(n_6628_o_0),
    .B(n_6630_o_0),
    .Y(n_6670_o_0));
 NAND2xp33_ASAP7_75t_R n_6671 (.A(n_6588_o_0),
    .B(n_6614_o_0),
    .Y(n_6671_o_0));
 AOI22xp33_ASAP7_75t_R n_6672 (.A1(n_6670_o_0),
    .A2(n_6624_o_0),
    .B1(n_6666_o_0),
    .B2(n_6671_o_0),
    .Y(n_6672_o_0));
 OA21x2_ASAP7_75t_R n_6673 (.A1(_00944_),
    .A2(n_6572_o_0),
    .B(n_6648_o_0),
    .Y(n_6673_o_0));
 XNOR2xp5_ASAP7_75t_R n_6674 (.A(_00946_),
    .B(n_6655_o_0),
    .Y(n_6674_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6675 (.A1(n_6669_o_0),
    .A2(n_6672_o_0),
    .B(n_6673_o_0),
    .C(n_6674_o_0),
    .Y(n_6675_o_0));
 OAI21xp33_ASAP7_75t_R n_6676 (.A1(n_6659_o_0),
    .A2(n_6668_o_0),
    .B(n_6675_o_0),
    .Y(n_6676_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6677 (.A1(n_6627_o_0),
    .A2(n_6635_o_0),
    .B(n_6658_o_0),
    .C(n_6676_o_0),
    .Y(n_6677_o_0));
 NOR2xp33_ASAP7_75t_R n_6678 (.A(n_6566_o_0),
    .B(n_6677_o_0),
    .Y(n_6678_o_0));
 INVx1_ASAP7_75t_R n_6679 (.A(n_6674_o_0),
    .Y(n_6679_o_0));
 AOI21xp33_ASAP7_75t_R n_6680 (.A1(n_6597_o_0),
    .A2(n_6598_o_0),
    .B(net2),
    .Y(n_6680_o_0));
 INVx1_ASAP7_75t_R n_6681 (.A(_00941_),
    .Y(n_6681_o_0));
 NOR2xp33_ASAP7_75t_R n_6682 (.A(_00549_),
    .B(net),
    .Y(n_6682_o_0));
 NOR3xp33_ASAP7_75t_R n_6683 (.A(n_6680_o_0),
    .B(n_6681_o_0),
    .C(n_6682_o_0),
    .Y(n_6683_o_0));
 OAI21xp33_ASAP7_75t_R n_6684 (.A1(n_6600_o_0),
    .A2(n_6683_o_0),
    .B(n_6588_o_0),
    .Y(n_6684_o_0));
 NAND2xp33_ASAP7_75t_R n_6685 (.A(n_6614_o_0),
    .B(n_6684_o_0),
    .Y(n_6685_o_0));
 NAND3xp33_ASAP7_75t_R n_6686 (.A(n_6661_o_0),
    .B(n_6644_o_0),
    .C(n_6630_o_0),
    .Y(n_6686_o_0));
 AOI21xp33_ASAP7_75t_R n_6687 (.A1(n_6685_o_0),
    .A2(n_6686_o_0),
    .B(n_6624_o_0),
    .Y(n_6687_o_0));
 AOI21xp33_ASAP7_75t_R n_6688 (.A1(n_6624_o_0),
    .A2(n_6670_o_0),
    .B(n_6687_o_0),
    .Y(n_6688_o_0));
 OAI31xp33_ASAP7_75t_R n_6689 (.A1(n_6600_o_0),
    .A2(n_6683_o_0),
    .A3(n_6588_o_0),
    .B(n_6637_o_0),
    .Y(n_6689_o_0));
 AOI21xp33_ASAP7_75t_R n_6690 (.A1(n_6630_o_0),
    .A2(n_6601_o_0),
    .B(n_6633_o_0),
    .Y(n_6690_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6691 (.A1(n_6594_o_0),
    .A2(_00941_),
    .B(n_6600_o_0),
    .C(n_6603_o_0),
    .Y(n_6691_o_0));
 NOR2xp33_ASAP7_75t_R n_6692 (.A(n_6691_o_0),
    .B(n_6630_o_0),
    .Y(n_6692_o_0));
 NAND2xp33_ASAP7_75t_R n_6693 (.A(n_6664_o_0),
    .B(n_6624_o_0),
    .Y(n_6693_o_0));
 OAI21xp33_ASAP7_75t_R n_6694 (.A1(n_6692_o_0),
    .A2(n_6693_o_0),
    .B(n_6673_o_0),
    .Y(n_6694_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6695 (.A1(n_6630_o_0),
    .A2(n_6689_o_0),
    .B(n_6690_o_0),
    .C(n_6694_o_0),
    .Y(n_6695_o_0));
 AOI21xp33_ASAP7_75t_R n_6696 (.A1(n_6573_o_0),
    .A2(n_6688_o_0),
    .B(n_6695_o_0),
    .Y(n_6696_o_0));
 INVx1_ASAP7_75t_R n_6697 (.A(n_6657_o_0),
    .Y(n_6697_o_0));
 NAND3xp33_ASAP7_75t_R n_6698 (.A(n_6630_o_0),
    .B(n_6588_o_0),
    .C(n_6601_o_0),
    .Y(n_6698_o_0));
 NAND2xp33_ASAP7_75t_R n_6699 (.A(n_6614_o_0),
    .B(n_6691_o_0),
    .Y(n_6699_o_0));
 AOI31xp33_ASAP7_75t_R n_6700 (.A1(n_6624_o_0),
    .A2(n_6698_o_0),
    .A3(n_6699_o_0),
    .B(n_6649_o_0),
    .Y(n_6700_o_0));
 OAI31xp33_ASAP7_75t_R n_6701 (.A1(n_6684_o_0),
    .A2(net55),
    .A3(n_6633_o_0),
    .B(n_6700_o_0),
    .Y(n_6701_o_0));
 INVx1_ASAP7_75t_R n_6702 (.A(n_6701_o_0),
    .Y(n_6702_o_0));
 AOI31xp33_ASAP7_75t_R n_6703 (.A1(n_6628_o_0),
    .A2(n_6603_o_0),
    .A3(n_6614_o_0),
    .B(n_6633_o_0),
    .Y(n_6703_o_0));
 NOR3xp33_ASAP7_75t_R n_6704 (.A(n_6684_o_0),
    .B(n_6666_o_0),
    .C(net55),
    .Y(n_6704_o_0));
 AOI211xp5_ASAP7_75t_R n_6705 (.A1(n_6703_o_0),
    .A2(n_6698_o_0),
    .B(n_6704_o_0),
    .C(n_6673_o_0),
    .Y(n_6705_o_0));
 NAND2xp33_ASAP7_75t_R n_6706 (.A(_00947_),
    .B(n_6564_o_0),
    .Y(n_6706_o_0));
 OAI21xp33_ASAP7_75t_R n_6707 (.A1(_00947_),
    .A2(n_6564_o_0),
    .B(n_6706_o_0),
    .Y(n_6707_o_0));
 INVx1_ASAP7_75t_R n_6708 (.A(n_6707_o_0),
    .Y(n_6708_o_0));
 OAI31xp33_ASAP7_75t_R n_6709 (.A1(n_6697_o_0),
    .A2(n_6702_o_0),
    .A3(n_6705_o_0),
    .B(n_6708_o_0),
    .Y(n_6709_o_0));
 AOI21xp33_ASAP7_75t_R n_6710 (.A1(n_6679_o_0),
    .A2(n_6696_o_0),
    .B(n_6709_o_0),
    .Y(n_6710_o_0));
 AOI211xp5_ASAP7_75t_R n_6711 (.A1(_00941_),
    .A2(n_6594_o_0),
    .B(n_6603_o_0),
    .C(n_6600_o_0),
    .Y(n_6711_o_0));
 NAND3xp33_ASAP7_75t_R n_6712 (.A(n_6661_o_0),
    .B(n_6711_o_0),
    .C(n_6614_o_0),
    .Y(n_6712_o_0));
 INVx1_ASAP7_75t_R n_6713 (.A(n_6689_o_0),
    .Y(n_6713_o_0));
 OAI21xp33_ASAP7_75t_R n_6714 (.A1(net55),
    .A2(n_6713_o_0),
    .B(n_6633_o_0),
    .Y(n_6714_o_0));
 NOR3xp33_ASAP7_75t_R n_6715 (.A(n_6624_o_0),
    .B(n_6691_o_0),
    .C(n_6614_o_0),
    .Y(n_6715_o_0));
 INVx1_ASAP7_75t_R n_6716 (.A(n_6715_o_0),
    .Y(n_6716_o_0));
 AO21x1_ASAP7_75t_R n_6717 (.A1(n_6714_o_0),
    .A2(n_6716_o_0),
    .B(n_6659_o_0),
    .Y(n_6717_o_0));
 NOR2xp33_ASAP7_75t_R n_6718 (.A(n_6614_o_0),
    .B(n_6601_o_0),
    .Y(n_6718_o_0));
 NAND2xp33_ASAP7_75t_R n_6719 (.A(n_6666_o_0),
    .B(n_6663_o_0),
    .Y(n_6719_o_0));
 OAI21xp33_ASAP7_75t_R n_6720 (.A1(n_6588_o_0),
    .A2(n_6628_o_0),
    .B(n_6630_o_0),
    .Y(n_6720_o_0));
 AOI31xp33_ASAP7_75t_R n_6721 (.A1(n_6624_o_0),
    .A2(n_6720_o_0),
    .A3(n_6671_o_0),
    .B(n_6659_o_0),
    .Y(n_6721_o_0));
 OAI21xp33_ASAP7_75t_R n_6722 (.A1(n_6718_o_0),
    .A2(n_6719_o_0),
    .B(n_6721_o_0),
    .Y(n_6722_o_0));
 AOI31xp33_ASAP7_75t_R n_6723 (.A1(n_6628_o_0),
    .A2(net55),
    .A3(n_6666_o_0),
    .B(n_6649_o_0),
    .Y(n_6723_o_0));
 OAI31xp33_ASAP7_75t_R n_6724 (.A1(n_6684_o_0),
    .A2(net55),
    .A3(n_6633_o_0),
    .B(n_6723_o_0),
    .Y(n_6724_o_0));
 NAND3xp33_ASAP7_75t_R n_6725 (.A(n_6630_o_0),
    .B(n_6603_o_0),
    .C(n_6601_o_0),
    .Y(n_6725_o_0));
 AND4x1_ASAP7_75t_R n_6726 (.A(n_6725_o_0),
    .B(n_6671_o_0),
    .C(n_6659_o_0),
    .D(n_6624_o_0),
    .Y(n_6726_o_0));
 AOI31xp33_ASAP7_75t_R n_6727 (.A1(n_6707_o_0),
    .A2(n_6722_o_0),
    .A3(n_6724_o_0),
    .B(n_6726_o_0),
    .Y(n_6727_o_0));
 NAND2xp33_ASAP7_75t_R n_6728 (.A(_00945_),
    .B(n_6556_o_0),
    .Y(n_6728_o_0));
 OAI21xp33_ASAP7_75t_R n_6729 (.A1(_00945_),
    .A2(n_6556_o_0),
    .B(n_6728_o_0),
    .Y(n_6729_o_0));
 INVx1_ASAP7_75t_R n_6730 (.A(n_6729_o_0),
    .Y(n_6730_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6731 (.A1(n_6712_o_0),
    .A2(n_6717_o_0),
    .B(n_6565_o_0),
    .C(n_6727_o_0),
    .D(n_6730_o_0),
    .Y(n_6731_o_0));
 NOR2xp33_ASAP7_75t_R n_6732 (.A(n_6697_o_0),
    .B(n_6730_o_0),
    .Y(n_6732_o_0));
 AOI31xp33_ASAP7_75t_R n_6733 (.A1(n_6614_o_0),
    .A2(n_6661_o_0),
    .A3(n_6644_o_0),
    .B(n_6573_o_0),
    .Y(n_6733_o_0));
 INVx1_ASAP7_75t_R n_6734 (.A(n_6733_o_0),
    .Y(n_6734_o_0));
 NOR2xp33_ASAP7_75t_R n_6735 (.A(n_6603_o_0),
    .B(n_6614_o_0),
    .Y(n_6735_o_0));
 AOI21xp33_ASAP7_75t_R n_6736 (.A1(n_6601_o_0),
    .A2(n_6735_o_0),
    .B(n_6624_o_0),
    .Y(n_6736_o_0));
 OAI21xp33_ASAP7_75t_R n_6737 (.A1(n_6630_o_0),
    .A2(n_6711_o_0),
    .B(n_6736_o_0),
    .Y(n_6737_o_0));
 INVx1_ASAP7_75t_R n_6738 (.A(n_6737_o_0),
    .Y(n_6738_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6739 (.A1(n_6614_o_0),
    .A2(n_6644_o_0),
    .B(n_6615_o_0),
    .C(n_6666_o_0),
    .Y(n_6739_o_0));
 NAND2xp33_ASAP7_75t_R n_6740 (.A(n_6601_o_0),
    .B(n_6630_o_0),
    .Y(n_6740_o_0));
 OAI321xp33_ASAP7_75t_R n_6741 (.A1(n_6630_o_0),
    .A2(n_6689_o_0),
    .A3(n_6624_o_0),
    .B1(n_6666_o_0),
    .B2(n_6740_o_0),
    .C(n_6649_o_0),
    .Y(n_6741_o_0));
 OAI31xp33_ASAP7_75t_R n_6742 (.A1(n_6734_o_0),
    .A2(n_6738_o_0),
    .A3(n_6739_o_0),
    .B(n_6741_o_0),
    .Y(n_6742_o_0));
 AOI211xp5_ASAP7_75t_R n_6743 (.A1(_00941_),
    .A2(n_6594_o_0),
    .B(n_6588_o_0),
    .C(n_6600_o_0),
    .Y(n_6743_o_0));
 AOI21xp33_ASAP7_75t_R n_6744 (.A1(n_6643_o_0),
    .A2(n_6639_o_0),
    .B(n_6603_o_0),
    .Y(n_6744_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6745 (.A1(n_6743_o_0),
    .A2(n_6744_o_0),
    .B(n_6614_o_0),
    .C(n_6666_o_0),
    .Y(n_6745_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6746 (.A1(n_6628_o_0),
    .A2(net55),
    .B(n_6641_o_0),
    .C(n_6661_o_0),
    .D(n_6745_o_0),
    .Y(n_6746_o_0));
 NAND3xp33_ASAP7_75t_R n_6747 (.A(n_6684_o_0),
    .B(n_6666_o_0),
    .C(n_6630_o_0),
    .Y(n_6747_o_0));
 OAI21xp33_ASAP7_75t_R n_6748 (.A1(n_6743_o_0),
    .A2(n_6744_o_0),
    .B(n_6630_o_0),
    .Y(n_6748_o_0));
 AOI211xp5_ASAP7_75t_R n_6749 (.A1(n_6603_o_0),
    .A2(n_6628_o_0),
    .B(n_6633_o_0),
    .C(n_6630_o_0),
    .Y(n_6749_o_0));
 AOI31xp33_ASAP7_75t_R n_6750 (.A1(n_6624_o_0),
    .A2(n_6748_o_0),
    .A3(n_6645_o_0),
    .B(n_6749_o_0),
    .Y(n_6750_o_0));
 AOI21xp33_ASAP7_75t_R n_6751 (.A1(n_6747_o_0),
    .A2(n_6750_o_0),
    .B(n_6573_o_0),
    .Y(n_6751_o_0));
 AOI211xp5_ASAP7_75t_R n_6752 (.A1(n_6649_o_0),
    .A2(n_6746_o_0),
    .B(n_6751_o_0),
    .C(n_6566_o_0),
    .Y(n_6752_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6753 (.A1(n_6566_o_0),
    .A2(n_6742_o_0),
    .B(n_6752_o_0),
    .C(n_6674_o_0),
    .Y(n_6753_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6754 (.A1(n_6731_o_0),
    .A2(n_6697_o_0),
    .B(n_6732_o_0),
    .C(n_6753_o_0),
    .Y(n_6754_o_0));
 OAI31xp33_ASAP7_75t_R n_6755 (.A1(n_6558_o_0),
    .A2(n_6678_o_0),
    .A3(n_6710_o_0),
    .B(n_6754_o_0),
    .Y(n_6755_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6756 (.A1(n_6604_o_0),
    .A2(n_6610_o_0),
    .B(n_6613_o_0),
    .C(n_6603_o_0),
    .Y(n_6756_o_0));
 OAI22xp33_ASAP7_75t_R n_6757 (.A1(n_6628_o_0),
    .A2(n_6756_o_0),
    .B1(n_6630_o_0),
    .B2(n_6691_o_0),
    .Y(n_6757_o_0));
 OAI21xp33_ASAP7_75t_R n_6758 (.A1(n_6624_o_0),
    .A2(n_6757_o_0),
    .B(n_6659_o_0),
    .Y(n_6758_o_0));
 NOR2xp33_ASAP7_75t_R n_6759 (.A(n_6601_o_0),
    .B(n_6630_o_0),
    .Y(n_6759_o_0));
 NOR3xp33_ASAP7_75t_R n_6760 (.A(n_6759_o_0),
    .B(n_6557_o_0),
    .C(n_6666_o_0),
    .Y(n_6760_o_0));
 NOR2xp33_ASAP7_75t_R n_6761 (.A(n_6630_o_0),
    .B(n_6628_o_0),
    .Y(n_6761_o_0));
 INVx1_ASAP7_75t_R n_6762 (.A(n_6761_o_0),
    .Y(n_6762_o_0));
 AOI21xp33_ASAP7_75t_R n_6763 (.A1(n_6628_o_0),
    .A2(n_6614_o_0),
    .B(n_6661_o_0),
    .Y(n_6763_o_0));
 AO21x1_ASAP7_75t_R n_6764 (.A1(n_6763_o_0),
    .A2(n_6670_o_0),
    .B(n_6557_o_0),
    .Y(n_6764_o_0));
 AOI21xp33_ASAP7_75t_R n_6765 (.A1(n_6634_o_0),
    .A2(n_6762_o_0),
    .B(n_6764_o_0),
    .Y(n_6765_o_0));
 AOI21xp33_ASAP7_75t_R n_6766 (.A1(n_6601_o_0),
    .A2(n_6603_o_0),
    .B(n_6661_o_0),
    .Y(n_6766_o_0));
 NAND2xp33_ASAP7_75t_R n_6767 (.A(n_6630_o_0),
    .B(n_6766_o_0),
    .Y(n_6767_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6768 (.A1(n_6601_o_0),
    .A2(n_6614_o_0),
    .B(n_6603_o_0),
    .C(n_6666_o_0),
    .Y(n_6768_o_0));
 NAND3xp33_ASAP7_75t_R n_6769 (.A(n_6602_o_0),
    .B(n_6624_o_0),
    .C(net55),
    .Y(n_6769_o_0));
 AND4x1_ASAP7_75t_R n_6770 (.A(n_6767_o_0),
    .B(n_6768_o_0),
    .C(n_6769_o_0),
    .D(n_6730_o_0),
    .Y(n_6770_o_0));
 OAI21xp33_ASAP7_75t_R n_6771 (.A1(n_6765_o_0),
    .A2(n_6770_o_0),
    .B(n_6573_o_0),
    .Y(n_6771_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6772 (.A1(n_6758_o_0),
    .A2(n_6760_o_0),
    .B(n_6771_o_0),
    .C(n_6679_o_0),
    .Y(n_6772_o_0));
 NOR2xp33_ASAP7_75t_R n_6773 (.A(n_6614_o_0),
    .B(n_6644_o_0),
    .Y(n_6773_o_0));
 INVx1_ASAP7_75t_R n_6774 (.A(n_6773_o_0),
    .Y(n_6774_o_0));
 NAND3xp33_ASAP7_75t_R n_6775 (.A(n_6661_o_0),
    .B(net55),
    .C(n_6603_o_0),
    .Y(n_6775_o_0));
 OAI211xp5_ASAP7_75t_R n_6776 (.A1(n_6774_o_0),
    .A2(n_6666_o_0),
    .B(n_6686_o_0),
    .C(n_6775_o_0),
    .Y(n_6776_o_0));
 OAI31xp33_ASAP7_75t_R n_6777 (.A1(n_6666_o_0),
    .A2(n_6689_o_0),
    .A3(n_6630_o_0),
    .B(n_6557_o_0),
    .Y(n_6777_o_0));
 OAI21xp33_ASAP7_75t_R n_6778 (.A1(n_6628_o_0),
    .A2(n_6615_o_0),
    .B(n_6624_o_0),
    .Y(n_6778_o_0));
 NOR2xp33_ASAP7_75t_R n_6779 (.A(n_6614_o_0),
    .B(n_6689_o_0),
    .Y(n_6779_o_0));
 AOI31xp33_ASAP7_75t_R n_6780 (.A1(n_6666_o_0),
    .A2(n_6685_o_0),
    .A3(n_6720_o_0),
    .B(n_6557_o_0),
    .Y(n_6780_o_0));
 OAI21xp33_ASAP7_75t_R n_6781 (.A1(n_6778_o_0),
    .A2(n_6779_o_0),
    .B(n_6780_o_0),
    .Y(n_6781_o_0));
 OA21x2_ASAP7_75t_R n_6782 (.A1(n_6776_o_0),
    .A2(n_6777_o_0),
    .B(n_6781_o_0),
    .Y(n_6782_o_0));
 NAND2xp33_ASAP7_75t_R n_6783 (.A(n_6666_o_0),
    .B(n_6671_o_0),
    .Y(n_6783_o_0));
 INVx1_ASAP7_75t_R n_6784 (.A(n_6725_o_0),
    .Y(n_6784_o_0));
 OAI21xp33_ASAP7_75t_R n_6785 (.A1(n_6783_o_0),
    .A2(n_6784_o_0),
    .B(n_6558_o_0),
    .Y(n_6785_o_0));
 AOI21xp33_ASAP7_75t_R n_6786 (.A1(n_6624_o_0),
    .A2(n_6748_o_0),
    .B(n_6785_o_0),
    .Y(n_6786_o_0));
 AO21x1_ASAP7_75t_R n_6787 (.A1(n_6763_o_0),
    .A2(n_6670_o_0),
    .B(n_6729_o_0),
    .Y(n_6787_o_0));
 AOI21xp33_ASAP7_75t_R n_6788 (.A1(n_6634_o_0),
    .A2(n_6645_o_0),
    .B(n_6787_o_0),
    .Y(n_6788_o_0));
 NOR3xp33_ASAP7_75t_R n_6789 (.A(n_6786_o_0),
    .B(n_6788_o_0),
    .C(n_6573_o_0),
    .Y(n_6789_o_0));
 AOI211xp5_ASAP7_75t_R n_6790 (.A1(n_6782_o_0),
    .A2(n_6649_o_0),
    .B(n_6789_o_0),
    .C(n_6657_o_0),
    .Y(n_6790_o_0));
 OAI21xp33_ASAP7_75t_R n_6791 (.A1(n_6778_o_0),
    .A2(n_6779_o_0),
    .B(n_6730_o_0),
    .Y(n_6791_o_0));
 AOI31xp33_ASAP7_75t_R n_6792 (.A1(n_6661_o_0),
    .A2(n_6711_o_0),
    .A3(n_6630_o_0),
    .B(n_6791_o_0),
    .Y(n_6792_o_0));
 OAI211xp5_ASAP7_75t_R n_6793 (.A1(n_6689_o_0),
    .A2(n_6630_o_0),
    .B(n_6666_o_0),
    .C(n_6664_o_0),
    .Y(n_6793_o_0));
 OAI21xp33_ASAP7_75t_R n_6794 (.A1(n_6743_o_0),
    .A2(n_6735_o_0),
    .B(n_6624_o_0),
    .Y(n_6794_o_0));
 AND3x1_ASAP7_75t_R n_6795 (.A(n_6793_o_0),
    .B(n_6794_o_0),
    .C(n_6558_o_0),
    .Y(n_6795_o_0));
 NOR3xp33_ASAP7_75t_R n_6796 (.A(n_6628_o_0),
    .B(n_6630_o_0),
    .C(n_6603_o_0),
    .Y(n_6796_o_0));
 AOI211xp5_ASAP7_75t_R n_6797 (.A1(n_6630_o_0),
    .A2(n_6689_o_0),
    .B(n_6796_o_0),
    .C(n_6661_o_0),
    .Y(n_6797_o_0));
 AOI31xp33_ASAP7_75t_R n_6798 (.A1(n_6666_o_0),
    .A2(n_6615_o_0),
    .A3(n_6774_o_0),
    .B(n_6797_o_0),
    .Y(n_6798_o_0));
 INVx1_ASAP7_75t_R n_6799 (.A(n_6662_o_0),
    .Y(n_6799_o_0));
 INVx1_ASAP7_75t_R n_6800 (.A(n_6718_o_0),
    .Y(n_6800_o_0));
 AOI211xp5_ASAP7_75t_R n_6801 (.A1(n_6601_o_0),
    .A2(n_6603_o_0),
    .B(n_6633_o_0),
    .C(n_6614_o_0),
    .Y(n_6801_o_0));
 AOI31xp33_ASAP7_75t_R n_6802 (.A1(n_6624_o_0),
    .A2(n_6799_o_0),
    .A3(n_6800_o_0),
    .B(n_6801_o_0),
    .Y(n_6802_o_0));
 AOI21xp33_ASAP7_75t_R n_6803 (.A1(n_6730_o_0),
    .A2(n_6802_o_0),
    .B(n_6673_o_0),
    .Y(n_6803_o_0));
 OAI21xp33_ASAP7_75t_R n_6804 (.A1(n_6730_o_0),
    .A2(n_6798_o_0),
    .B(n_6803_o_0),
    .Y(n_6804_o_0));
 OAI31xp33_ASAP7_75t_R n_6805 (.A1(n_6573_o_0),
    .A2(n_6792_o_0),
    .A3(n_6795_o_0),
    .B(n_6804_o_0),
    .Y(n_6805_o_0));
 NOR2xp33_ASAP7_75t_R n_6806 (.A(n_6588_o_0),
    .B(n_6628_o_0),
    .Y(n_6806_o_0));
 OA21x2_ASAP7_75t_R n_6807 (.A1(net55),
    .A2(n_6806_o_0),
    .B(n_6745_o_0),
    .Y(n_6807_o_0));
 AOI31xp33_ASAP7_75t_R n_6808 (.A1(net55),
    .A2(n_6661_o_0),
    .A3(n_6711_o_0),
    .B(n_6673_o_0),
    .Y(n_6808_o_0));
 OAI211xp5_ASAP7_75t_R n_6809 (.A1(n_6761_o_0),
    .A2(n_6666_o_0),
    .B(n_6808_o_0),
    .C(n_6800_o_0),
    .Y(n_6809_o_0));
 OAI31xp33_ASAP7_75t_R n_6810 (.A1(n_6573_o_0),
    .A2(n_6738_o_0),
    .A3(n_6807_o_0),
    .B(n_6809_o_0),
    .Y(n_6810_o_0));
 INVx1_ASAP7_75t_R n_6811 (.A(n_6769_o_0),
    .Y(n_6811_o_0));
 AO21x1_ASAP7_75t_R n_6812 (.A1(n_6690_o_0),
    .A2(n_6629_o_0),
    .B(n_6649_o_0),
    .Y(n_6812_o_0));
 NAND2xp33_ASAP7_75t_R n_6813 (.A(n_6624_o_0),
    .B(n_6748_o_0),
    .Y(n_6813_o_0));
 AOI31xp33_ASAP7_75t_R n_6814 (.A1(n_6666_o_0),
    .A2(n_6670_o_0),
    .A3(n_6615_o_0),
    .B(n_6659_o_0),
    .Y(n_6814_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6815 (.A1(net55),
    .A2(n_6588_o_0),
    .B(n_6813_o_0),
    .C(n_6814_o_0),
    .Y(n_6815_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6816 (.A1(n_6811_o_0),
    .A2(n_6812_o_0),
    .B(n_6815_o_0),
    .C(n_6729_o_0),
    .Y(n_6816_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6817 (.A1(n_6810_o_0),
    .A2(n_6729_o_0),
    .B(n_6816_o_0),
    .C(n_6657_o_0),
    .Y(n_6817_o_0));
 OAI211xp5_ASAP7_75t_R n_6818 (.A1(n_6805_o_0),
    .A2(n_6657_o_0),
    .B(n_6566_o_0),
    .C(n_6817_o_0),
    .Y(n_6818_o_0));
 OAI31xp33_ASAP7_75t_R n_6819 (.A1(n_6708_o_0),
    .A2(n_6772_o_0),
    .A3(n_6790_o_0),
    .B(n_6818_o_0),
    .Y(n_6819_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6820 (.A1(n_6588_o_0),
    .A2(n_6630_o_0),
    .B(n_6601_o_0),
    .C(n_6661_o_0),
    .Y(n_6820_o_0));
 AOI31xp33_ASAP7_75t_R n_6821 (.A1(n_6666_o_0),
    .A2(n_6799_o_0),
    .A3(n_6670_o_0),
    .B(n_6820_o_0),
    .Y(n_6821_o_0));
 OAI21xp33_ASAP7_75t_R n_6822 (.A1(n_6673_o_0),
    .A2(n_6821_o_0),
    .B(n_6558_o_0),
    .Y(n_6822_o_0));
 INVx1_ASAP7_75t_R n_6823 (.A(n_6690_o_0),
    .Y(n_6823_o_0));
 NOR2xp33_ASAP7_75t_R n_6824 (.A(n_6630_o_0),
    .B(n_6689_o_0),
    .Y(n_6824_o_0));
 INVx1_ASAP7_75t_R n_6825 (.A(n_6664_o_0),
    .Y(n_6825_o_0));
 NOR2xp33_ASAP7_75t_R n_6826 (.A(n_6630_o_0),
    .B(n_6711_o_0),
    .Y(n_6826_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6827 (.A1(n_6825_o_0),
    .A2(n_6601_o_0),
    .B(n_6826_o_0),
    .C(n_6633_o_0),
    .Y(n_6827_o_0));
 OA211x2_ASAP7_75t_R n_6828 (.A1(n_6823_o_0),
    .A2(n_6824_o_0),
    .B(n_6827_o_0),
    .C(n_6659_o_0),
    .Y(n_6828_o_0));
 OAI21xp33_ASAP7_75t_R n_6829 (.A1(n_6822_o_0),
    .A2(n_6828_o_0),
    .B(n_6565_o_0),
    .Y(n_6829_o_0));
 NAND2xp33_ASAP7_75t_R n_6830 (.A(n_6558_o_0),
    .B(n_6829_o_0),
    .Y(n_6830_o_0));
 OAI21xp33_ASAP7_75t_R n_6831 (.A1(n_6600_o_0),
    .A2(n_6683_o_0),
    .B(n_6630_o_0),
    .Y(n_6831_o_0));
 AOI321xp33_ASAP7_75t_R n_6832 (.A1(n_6630_o_0),
    .A2(n_6640_o_0),
    .A3(n_6637_o_0),
    .B1(n_6831_o_0),
    .B2(n_6628_o_0),
    .C(n_6633_o_0),
    .Y(n_6832_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6833 (.A1(n_6756_o_0),
    .A2(n_6624_o_0),
    .B(n_6832_o_0),
    .C(n_6645_o_0),
    .Y(n_6833_o_0));
 INVx1_ASAP7_75t_R n_6834 (.A(n_6720_o_0),
    .Y(n_6834_o_0));
 OAI211xp5_ASAP7_75t_R n_6835 (.A1(n_6834_o_0),
    .A2(n_6778_o_0),
    .B(n_6719_o_0),
    .C(n_6673_o_0),
    .Y(n_6835_o_0));
 OAI21xp33_ASAP7_75t_R n_6836 (.A1(n_6673_o_0),
    .A2(n_6833_o_0),
    .B(n_6835_o_0),
    .Y(n_6836_o_0));
 OAI21xp33_ASAP7_75t_R n_6837 (.A1(n_6836_o_0),
    .A2(n_6829_o_0),
    .B(n_6557_o_0),
    .Y(n_6837_o_0));
 NOR2xp33_ASAP7_75t_R n_6838 (.A(n_6588_o_0),
    .B(n_6614_o_0),
    .Y(n_6838_o_0));
 OAI21xp33_ASAP7_75t_R n_6839 (.A1(n_6838_o_0),
    .A2(n_6778_o_0),
    .B(n_6573_o_0),
    .Y(n_6839_o_0));
 AOI21xp33_ASAP7_75t_R n_6840 (.A1(n_6703_o_0),
    .A2(n_6725_o_0),
    .B(n_6839_o_0),
    .Y(n_6840_o_0));
 INVx1_ASAP7_75t_R n_6841 (.A(n_6826_o_0),
    .Y(n_6841_o_0));
 OAI31xp33_ASAP7_75t_R n_6842 (.A1(n_6633_o_0),
    .A2(net55),
    .A3(n_6644_o_0),
    .B(n_6673_o_0),
    .Y(n_6842_o_0));
 AOI31xp33_ASAP7_75t_R n_6843 (.A1(n_6624_o_0),
    .A2(n_6748_o_0),
    .A3(n_6841_o_0),
    .B(n_6842_o_0),
    .Y(n_6843_o_0));
 NOR3xp33_ASAP7_75t_R n_6844 (.A(n_6624_o_0),
    .B(n_6630_o_0),
    .C(n_6628_o_0),
    .Y(n_6844_o_0));
 AOI22xp33_ASAP7_75t_R n_6845 (.A1(n_6663_o_0),
    .A2(n_6666_o_0),
    .B1(n_6740_o_0),
    .B2(n_6624_o_0),
    .Y(n_6845_o_0));
 AOI21xp33_ASAP7_75t_R n_6846 (.A1(n_6673_o_0),
    .A2(n_6845_o_0),
    .B(n_6730_o_0),
    .Y(n_6846_o_0));
 OAI31xp33_ASAP7_75t_R n_6847 (.A1(n_6820_o_0),
    .A2(n_6844_o_0),
    .A3(n_6659_o_0),
    .B(n_6846_o_0),
    .Y(n_6847_o_0));
 OAI31xp33_ASAP7_75t_R n_6848 (.A1(n_6558_o_0),
    .A2(n_6840_o_0),
    .A3(n_6843_o_0),
    .B(n_6847_o_0),
    .Y(n_6848_o_0));
 AOI21xp33_ASAP7_75t_R n_6849 (.A1(n_6566_o_0),
    .A2(n_6848_o_0),
    .B(n_6679_o_0),
    .Y(n_6849_o_0));
 AO21x1_ASAP7_75t_R n_6850 (.A1(n_6557_o_0),
    .A2(n_6836_o_0),
    .B(n_6829_o_0),
    .Y(n_6850_o_0));
 OAI21xp33_ASAP7_75t_R n_6851 (.A1(n_6743_o_0),
    .A2(n_6744_o_0),
    .B(n_6614_o_0),
    .Y(n_6851_o_0));
 AOI21xp33_ASAP7_75t_R n_6852 (.A1(n_6646_o_0),
    .A2(n_6851_o_0),
    .B(n_6666_o_0),
    .Y(n_6852_o_0));
 AOI21xp33_ASAP7_75t_R n_6853 (.A1(n_6690_o_0),
    .A2(n_6685_o_0),
    .B(n_6852_o_0),
    .Y(n_6853_o_0));
 AOI21xp33_ASAP7_75t_R n_6854 (.A1(n_6628_o_0),
    .A2(n_6588_o_0),
    .B(n_6661_o_0),
    .Y(n_6854_o_0));
 HAxp5_ASAP7_75t_R n_6855 (.A(n_6630_o_0),
    .B(n_6601_o_0),
    .CON(n_6855_o_0),
    .SN(n_6855_o_1));
 AOI21xp33_ASAP7_75t_R n_6856 (.A1(n_6854_o_0),
    .A2(n_6855_o_0),
    .B(n_6649_o_0),
    .Y(n_6856_o_0));
 INVx1_ASAP7_75t_R n_6857 (.A(n_6856_o_0),
    .Y(n_6857_o_0));
 OAI21xp33_ASAP7_75t_R n_6858 (.A1(n_6673_o_0),
    .A2(n_6853_o_0),
    .B(n_6857_o_0),
    .Y(n_6858_o_0));
 OAI311xp33_ASAP7_75t_R n_6859 (.A1(n_6624_o_0),
    .A2(n_6649_o_0),
    .A3(n_6759_o_0),
    .B1(n_6729_o_0),
    .C1(n_6858_o_0),
    .Y(n_6859_o_0));
 OAI21xp33_ASAP7_75t_R n_6860 (.A1(n_6630_o_0),
    .A2(n_6689_o_0),
    .B(n_6690_o_0),
    .Y(n_6860_o_0));
 NAND2xp33_ASAP7_75t_R n_6861 (.A(n_6664_o_0),
    .B(n_6763_o_0),
    .Y(n_6861_o_0));
 NAND2xp33_ASAP7_75t_R n_6862 (.A(n_6588_o_0),
    .B(n_6601_o_0),
    .Y(n_6862_o_0));
 OAI21xp33_ASAP7_75t_R n_6863 (.A1(n_6624_o_0),
    .A2(n_6740_o_0),
    .B(n_6659_o_0),
    .Y(n_6863_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6864 (.A1(n_6862_o_0),
    .A2(net55),
    .B(n_6745_o_0),
    .C(n_6863_o_0),
    .Y(n_6864_o_0));
 AOI31xp33_ASAP7_75t_R n_6865 (.A1(n_6649_o_0),
    .A2(n_6860_o_0),
    .A3(n_6861_o_0),
    .B(n_6864_o_0),
    .Y(n_6865_o_0));
 OAI211xp5_ASAP7_75t_R n_6866 (.A1(n_6865_o_0),
    .A2(n_6558_o_0),
    .B(n_6679_o_0),
    .C(n_6708_o_0),
    .Y(n_6866_o_0));
 INVx1_ASAP7_75t_R n_6867 (.A(n_6860_o_0),
    .Y(n_6867_o_0));
 INVx1_ASAP7_75t_R n_6868 (.A(n_6861_o_0),
    .Y(n_6868_o_0));
 OAI21xp33_ASAP7_75t_R n_6869 (.A1(n_6862_o_0),
    .A2(n_6614_o_0),
    .B(n_6745_o_0),
    .Y(n_6869_o_0));
 OAI211xp5_ASAP7_75t_R n_6870 (.A1(n_6624_o_0),
    .A2(n_6740_o_0),
    .B(n_6869_o_0),
    .C(n_6659_o_0),
    .Y(n_6870_o_0));
 OAI31xp33_ASAP7_75t_R n_6871 (.A1(n_6673_o_0),
    .A2(n_6867_o_0),
    .A3(n_6868_o_0),
    .B(n_6870_o_0),
    .Y(n_6871_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6872 (.A1(n_6871_o_0),
    .A2(n_6557_o_0),
    .B(n_6707_o_0),
    .C(n_6679_o_0),
    .Y(n_6872_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6873 (.A1(n_6630_o_0),
    .A2(n_6691_o_0),
    .B(n_6634_o_0),
    .C(n_6649_o_0),
    .Y(n_6873_o_0));
 OAI21xp33_ASAP7_75t_R n_6874 (.A1(n_6689_o_0),
    .A2(net55),
    .B(n_6745_o_0),
    .Y(n_6874_o_0));
 OAI31xp33_ASAP7_75t_R n_6875 (.A1(n_6628_o_0),
    .A2(n_6588_o_0),
    .A3(n_6630_o_0),
    .B(n_6666_o_0),
    .Y(n_6875_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6876 (.A1(n_6630_o_0),
    .A2(n_6603_o_0),
    .B(n_6875_o_0),
    .C(n_6573_o_0),
    .Y(n_6876_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6877 (.A1(n_6646_o_0),
    .A2(n_6763_o_0),
    .B(n_6876_o_0),
    .C(n_6557_o_0),
    .Y(n_6877_o_0));
 AOI21xp33_ASAP7_75t_R n_6878 (.A1(n_6630_o_0),
    .A2(n_6603_o_0),
    .B(n_6796_o_0),
    .Y(n_6878_o_0));
 AOI21xp33_ASAP7_75t_R n_6879 (.A1(n_6573_o_0),
    .A2(n_6875_o_0),
    .B(n_6715_o_0),
    .Y(n_6879_o_0));
 OAI21xp33_ASAP7_75t_R n_6880 (.A1(n_6603_o_0),
    .A2(n_6628_o_0),
    .B(net55),
    .Y(n_6880_o_0));
 OAI21xp33_ASAP7_75t_R n_6881 (.A1(n_6628_o_0),
    .A2(n_6666_o_0),
    .B(n_6630_o_0),
    .Y(n_6881_o_0));
 AOI31xp33_ASAP7_75t_R n_6882 (.A1(n_6880_o_0),
    .A2(n_6881_o_0),
    .A3(n_6673_o_0),
    .B(n_6730_o_0),
    .Y(n_6882_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6883 (.A1(n_6878_o_0),
    .A2(n_6624_o_0),
    .B(n_6879_o_0),
    .C(n_6882_o_0),
    .Y(n_6883_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6884 (.A1(n_6873_o_0),
    .A2(n_6874_o_0),
    .B(n_6877_o_0),
    .C(n_6883_o_0),
    .Y(n_6884_o_0));
 NOR2xp33_ASAP7_75t_R n_6885 (.A(n_6566_o_0),
    .B(n_6884_o_0),
    .Y(n_6885_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6886 (.A1(n_6859_o_0),
    .A2(n_6866_o_0),
    .B(n_6872_o_0),
    .C(n_6885_o_0),
    .Y(n_6886_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6887 (.A1(n_6830_o_0),
    .A2(n_6837_o_0),
    .B(n_6849_o_0),
    .C(n_6850_o_0),
    .D(n_6886_o_0),
    .Y(n_6887_o_0));
 AOI211xp5_ASAP7_75t_R n_6888 (.A1(net55),
    .A2(n_6628_o_0),
    .B(n_6735_o_0),
    .C(n_6624_o_0),
    .Y(n_6888_o_0));
 OAI31xp33_ASAP7_75t_R n_6889 (.A1(n_6673_o_0),
    .A2(n_6888_o_0),
    .A3(n_6745_o_0),
    .B(n_6674_o_0),
    .Y(n_6889_o_0));
 OAI21xp33_ASAP7_75t_R n_6890 (.A1(n_6601_o_0),
    .A2(n_6630_o_0),
    .B(n_6624_o_0),
    .Y(n_6890_o_0));
 OAI21xp33_ASAP7_75t_R n_6891 (.A1(n_6890_o_0),
    .A2(n_6641_o_0),
    .B(n_6673_o_0),
    .Y(n_6891_o_0));
 AOI21xp33_ASAP7_75t_R n_6892 (.A1(n_6634_o_0),
    .A2(n_6602_o_0),
    .B(n_6891_o_0),
    .Y(n_6892_o_0));
 OAI311xp33_ASAP7_75t_R n_6893 (.A1(net55),
    .A2(n_6744_o_0),
    .A3(n_6743_o_0),
    .B1(n_6666_o_0),
    .C1(n_6699_o_0),
    .Y(n_6893_o_0));
 OAI31xp33_ASAP7_75t_R n_6894 (.A1(n_6661_o_0),
    .A2(n_6662_o_0),
    .A3(n_6718_o_0),
    .B(n_6893_o_0),
    .Y(n_6894_o_0));
 AOI31xp33_ASAP7_75t_R n_6895 (.A1(n_6666_o_0),
    .A2(n_6756_o_0),
    .A3(n_6602_o_0),
    .B(n_6649_o_0),
    .Y(n_6895_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6896 (.A1(n_6661_o_0),
    .A2(n_6669_o_0),
    .B(n_6895_o_0),
    .C(n_6674_o_0),
    .Y(n_6896_o_0));
 OAI21xp33_ASAP7_75t_R n_6897 (.A1(n_6659_o_0),
    .A2(n_6894_o_0),
    .B(n_6896_o_0),
    .Y(n_6897_o_0));
 OA21x2_ASAP7_75t_R n_6898 (.A1(n_6889_o_0),
    .A2(n_6892_o_0),
    .B(n_6897_o_0),
    .Y(n_6898_o_0));
 AOI21xp33_ASAP7_75t_R n_6899 (.A1(n_6630_o_0),
    .A2(n_6689_o_0),
    .B(n_6624_o_0),
    .Y(n_6899_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6900 (.A1(n_6603_o_0),
    .A2(n_6628_o_0),
    .B(n_6630_o_0),
    .C(n_6899_o_0),
    .Y(n_6900_o_0));
 INVx1_ASAP7_75t_R n_6901 (.A(n_6900_o_0),
    .Y(n_6901_o_0));
 OAI21xp33_ASAP7_75t_R n_6902 (.A1(n_6614_o_0),
    .A2(n_6691_o_0),
    .B(n_6671_o_0),
    .Y(n_6902_o_0));
 AOI21xp33_ASAP7_75t_R n_6903 (.A1(n_6763_o_0),
    .A2(n_6902_o_0),
    .B(n_6649_o_0),
    .Y(n_6903_o_0));
 OAI21xp33_ASAP7_75t_R n_6904 (.A1(n_6793_o_0),
    .A2(n_6718_o_0),
    .B(n_6903_o_0),
    .Y(n_6904_o_0));
 OAI21xp33_ASAP7_75t_R n_6905 (.A1(n_6626_o_0),
    .A2(n_6901_o_0),
    .B(n_6904_o_0),
    .Y(n_6905_o_0));
 NAND2xp33_ASAP7_75t_R n_6906 (.A(n_6661_o_0),
    .B(n_6832_o_0),
    .Y(n_6906_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6907 (.A1(n_6841_o_0),
    .A2(n_6720_o_0),
    .B(n_6832_o_0),
    .C(n_6624_o_0),
    .Y(n_6907_o_0));
 AO21x1_ASAP7_75t_R n_6908 (.A1(n_6646_o_0),
    .A2(n_6671_o_0),
    .B(n_6624_o_0),
    .Y(n_6908_o_0));
 NAND2xp33_ASAP7_75t_R n_6909 (.A(n_6630_o_0),
    .B(n_6684_o_0),
    .Y(n_6909_o_0));
 AOI21xp33_ASAP7_75t_R n_6910 (.A1(n_6909_o_0),
    .A2(n_6745_o_0),
    .B(n_6673_o_0),
    .Y(n_6910_o_0));
 AOI21xp33_ASAP7_75t_R n_6911 (.A1(n_6908_o_0),
    .A2(n_6910_o_0),
    .B(n_6679_o_0),
    .Y(n_6911_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6912 (.A1(n_6906_o_0),
    .A2(n_6907_o_0),
    .B(n_6573_o_0),
    .C(n_6911_o_0),
    .D(n_6558_o_0),
    .Y(n_6912_o_0));
 OAI21xp33_ASAP7_75t_R n_6913 (.A1(n_6657_o_0),
    .A2(n_6905_o_0),
    .B(n_6912_o_0),
    .Y(n_6913_o_0));
 OAI21xp33_ASAP7_75t_R n_6914 (.A1(n_6730_o_0),
    .A2(n_6898_o_0),
    .B(n_6913_o_0),
    .Y(n_6914_o_0));
 AOI21xp33_ASAP7_75t_R n_6915 (.A1(n_6671_o_0),
    .A2(n_6646_o_0),
    .B(n_6666_o_0),
    .Y(n_6915_o_0));
 INVx1_ASAP7_75t_R n_6916 (.A(n_6915_o_0),
    .Y(n_6916_o_0));
 OAI21xp33_ASAP7_75t_R n_6917 (.A1(n_6630_o_0),
    .A2(n_6806_o_0),
    .B(n_6899_o_0),
    .Y(n_6917_o_0));
 AOI211xp5_ASAP7_75t_R n_6918 (.A1(n_6690_o_0),
    .A2(n_6629_o_0),
    .B(n_6739_o_0),
    .C(n_6649_o_0),
    .Y(n_6918_o_0));
 AOI31xp33_ASAP7_75t_R n_6919 (.A1(n_6649_o_0),
    .A2(n_6916_o_0),
    .A3(n_6917_o_0),
    .B(n_6918_o_0),
    .Y(n_6919_o_0));
 OAI21xp33_ASAP7_75t_R n_6920 (.A1(n_6614_o_0),
    .A2(n_6691_o_0),
    .B(n_6624_o_0),
    .Y(n_6920_o_0));
 INVx1_ASAP7_75t_R n_6921 (.A(n_6920_o_0),
    .Y(n_6921_o_0));
 INVx1_ASAP7_75t_R n_6922 (.A(n_6873_o_0),
    .Y(n_6922_o_0));
 AOI211xp5_ASAP7_75t_R n_6923 (.A1(n_6640_o_0),
    .A2(n_6637_o_0),
    .B(n_6624_o_0),
    .C(n_6614_o_0),
    .Y(n_6923_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6924 (.A1(n_6923_o_0),
    .A2(n_6704_o_0),
    .B(n_6573_o_0),
    .C(n_6697_o_0),
    .Y(n_6924_o_0));
 OAI21xp33_ASAP7_75t_R n_6925 (.A1(n_6921_o_0),
    .A2(n_6922_o_0),
    .B(n_6924_o_0),
    .Y(n_6925_o_0));
 OAI21xp33_ASAP7_75t_R n_6926 (.A1(n_6674_o_0),
    .A2(n_6919_o_0),
    .B(n_6925_o_0),
    .Y(n_6926_o_0));
 OAI21xp33_ASAP7_75t_R n_6927 (.A1(n_6603_o_0),
    .A2(n_6666_o_0),
    .B(n_6630_o_0),
    .Y(n_6927_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6928 (.A1(n_6806_o_0),
    .A2(n_6633_o_0),
    .B(n_6630_o_0),
    .C(n_6927_o_0),
    .Y(n_6928_o_0));
 OAI21xp33_ASAP7_75t_R n_6929 (.A1(n_6630_o_0),
    .A2(n_6603_o_0),
    .B(n_6899_o_0),
    .Y(n_6929_o_0));
 AOI21xp33_ASAP7_75t_R n_6930 (.A1(n_6637_o_0),
    .A2(n_6640_o_0),
    .B(n_6630_o_0),
    .Y(n_6930_o_0));
 OAI31xp33_ASAP7_75t_R n_6931 (.A1(net55),
    .A2(n_6684_o_0),
    .A3(n_6666_o_0),
    .B(n_6649_o_0),
    .Y(n_6931_o_0));
 AOI221xp5_ASAP7_75t_R n_6932 (.A1(n_6633_o_0),
    .A2(n_6930_o_0),
    .B1(n_6703_o_0),
    .B2(n_6855_o_0),
    .C(n_6931_o_0),
    .Y(n_6932_o_0));
 AOI31xp33_ASAP7_75t_R n_6933 (.A1(n_6659_o_0),
    .A2(n_6928_o_0),
    .A3(n_6929_o_0),
    .B(n_6932_o_0),
    .Y(n_6933_o_0));
 AOI21xp33_ASAP7_75t_R n_6934 (.A1(n_6630_o_0),
    .A2(n_6603_o_0),
    .B(n_6875_o_0),
    .Y(n_6934_o_0));
 OAI21xp33_ASAP7_75t_R n_6935 (.A1(n_6691_o_0),
    .A2(n_6666_o_0),
    .B(net55),
    .Y(n_6935_o_0));
 OAI21xp33_ASAP7_75t_R n_6936 (.A1(n_6603_o_0),
    .A2(n_6666_o_0),
    .B(n_6630_o_0),
    .Y(n_6936_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6937 (.A1(n_6935_o_0),
    .A2(n_6936_o_0),
    .B(n_6758_o_0),
    .C(n_6697_o_0),
    .Y(n_6937_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6938 (.A1(n_6649_o_0),
    .A2(n_6934_o_0),
    .B(n_6937_o_0),
    .C(n_6729_o_0),
    .Y(n_6938_o_0));
 AOI21xp33_ASAP7_75t_R n_6939 (.A1(n_6674_o_0),
    .A2(n_6933_o_0),
    .B(n_6938_o_0),
    .Y(n_6939_o_0));
 AOI211xp5_ASAP7_75t_R n_6940 (.A1(n_6926_o_0),
    .A2(n_6557_o_0),
    .B(n_6566_o_0),
    .C(n_6939_o_0),
    .Y(n_6940_o_0));
 AO21x1_ASAP7_75t_R n_6941 (.A1(n_6914_o_0),
    .A2(n_6566_o_0),
    .B(n_6940_o_0),
    .Y(n_6941_o_0));
 AOI32xp33_ASAP7_75t_R n_6942 (.A1(n_6666_o_0),
    .A2(n_6799_o_0),
    .A3(n_6670_o_0),
    .B1(n_6698_o_0),
    .B2(n_6763_o_0),
    .Y(n_6942_o_0));
 OAI21xp33_ASAP7_75t_R n_6943 (.A1(n_6666_o_0),
    .A2(n_6774_o_0),
    .B(n_6659_o_0),
    .Y(n_6943_o_0));
 OAI21xp33_ASAP7_75t_R n_6944 (.A1(n_6666_o_0),
    .A2(n_6762_o_0),
    .B(n_6737_o_0),
    .Y(n_6944_o_0));
 OAI21xp33_ASAP7_75t_R n_6945 (.A1(n_6943_o_0),
    .A2(n_6944_o_0),
    .B(n_6558_o_0),
    .Y(n_6945_o_0));
 AOI21xp33_ASAP7_75t_R n_6946 (.A1(n_6649_o_0),
    .A2(n_6942_o_0),
    .B(n_6945_o_0),
    .Y(n_6946_o_0));
 OAI311xp33_ASAP7_75t_R n_6947 (.A1(n_6666_o_0),
    .A2(n_6630_o_0),
    .A3(n_6689_o_0),
    .B1(n_6646_o_0),
    .C1(n_6712_o_0),
    .Y(n_6947_o_0));
 INVx1_ASAP7_75t_R n_6948 (.A(n_6947_o_0),
    .Y(n_6948_o_0));
 NAND2xp33_ASAP7_75t_R n_6949 (.A(n_6666_o_0),
    .B(n_6720_o_0),
    .Y(n_6949_o_0));
 OAI21xp33_ASAP7_75t_R n_6950 (.A1(n_6930_o_0),
    .A2(n_6949_o_0),
    .B(n_6673_o_0),
    .Y(n_6950_o_0));
 AOI31xp33_ASAP7_75t_R n_6951 (.A1(n_6624_o_0),
    .A2(n_6699_o_0),
    .A3(n_6698_o_0),
    .B(n_6950_o_0),
    .Y(n_6951_o_0));
 AOI211xp5_ASAP7_75t_R n_6952 (.A1(n_6649_o_0),
    .A2(n_6948_o_0),
    .B(n_6951_o_0),
    .C(n_6729_o_0),
    .Y(n_6952_o_0));
 AOI21xp33_ASAP7_75t_R n_6953 (.A1(n_6614_o_0),
    .A2(n_6691_o_0),
    .B(n_6666_o_0),
    .Y(n_6953_o_0));
 AOI211xp5_ASAP7_75t_R n_6954 (.A1(n_6630_o_0),
    .A2(n_6644_o_0),
    .B(n_6953_o_0),
    .C(n_6673_o_0),
    .Y(n_6954_o_0));
 OA211x2_ASAP7_75t_R n_6955 (.A1(n_6693_o_0),
    .A2(n_6761_o_0),
    .B(n_6768_o_0),
    .C(n_6673_o_0),
    .Y(n_6955_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6956 (.A1(n_6588_o_0),
    .A2(n_6630_o_0),
    .B(n_6628_o_0),
    .C(n_6661_o_0),
    .Y(n_6956_o_0));
 AOI211xp5_ASAP7_75t_R n_6957 (.A1(n_6628_o_0),
    .A2(n_6630_o_0),
    .B(n_6624_o_0),
    .C(n_6743_o_0),
    .Y(n_6957_o_0));
 NAND2xp33_ASAP7_75t_R n_6958 (.A(n_6614_o_0),
    .B(n_6628_o_0),
    .Y(n_6958_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6959 (.A1(n_6664_o_0),
    .A2(n_6958_o_0),
    .B(n_6624_o_0),
    .C(n_6856_o_0),
    .Y(n_6959_o_0));
 OAI31xp33_ASAP7_75t_R n_6960 (.A1(n_6673_o_0),
    .A2(n_6956_o_0),
    .A3(n_6957_o_0),
    .B(n_6959_o_0),
    .Y(n_6960_o_0));
 OAI321xp33_ASAP7_75t_R n_6961 (.A1(n_6729_o_0),
    .A2(n_6954_o_0),
    .A3(n_6955_o_0),
    .B1(n_6960_o_0),
    .B2(n_6557_o_0),
    .C(n_6679_o_0),
    .Y(n_6961_o_0));
 OAI31xp33_ASAP7_75t_R n_6962 (.A1(n_6946_o_0),
    .A2(n_6952_o_0),
    .A3(n_6697_o_0),
    .B(n_6961_o_0),
    .Y(n_6962_o_0));
 OAI21xp33_ASAP7_75t_R n_6963 (.A1(n_6614_o_0),
    .A2(n_6711_o_0),
    .B(n_6666_o_0),
    .Y(n_6963_o_0));
 OAI21xp33_ASAP7_75t_R n_6964 (.A1(n_6963_o_0),
    .A2(n_6824_o_0),
    .B(n_6730_o_0),
    .Y(n_6964_o_0));
 AOI31xp33_ASAP7_75t_R n_6965 (.A1(n_6624_o_0),
    .A2(n_6671_o_0),
    .A3(n_6725_o_0),
    .B(n_6964_o_0),
    .Y(n_6965_o_0));
 OAI21xp33_ASAP7_75t_R n_6966 (.A1(n_6603_o_0),
    .A2(n_6633_o_0),
    .B(n_6630_o_0),
    .Y(n_6966_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6967 (.A1(n_6624_o_0),
    .A2(n_6799_o_0),
    .B(n_6966_o_0),
    .C(n_6557_o_0),
    .Y(n_6967_o_0));
 INVx1_ASAP7_75t_R n_6968 (.A(n_6778_o_0),
    .Y(n_6968_o_0));
 AOI21xp33_ASAP7_75t_R n_6969 (.A1(n_6614_o_0),
    .A2(n_6684_o_0),
    .B(n_6633_o_0),
    .Y(n_6969_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_6970 (.A1(n_6601_o_0),
    .A2(n_6630_o_0),
    .B(n_6747_o_0),
    .C(n_6633_o_0),
    .Y(n_6970_o_0));
 OAI321xp33_ASAP7_75t_R n_6971 (.A1(n_6729_o_0),
    .A2(n_6968_o_0),
    .A3(n_6969_o_0),
    .B1(n_6764_o_0),
    .B2(n_6970_o_0),
    .C(n_6649_o_0),
    .Y(n_6971_o_0));
 OAI31xp33_ASAP7_75t_R n_6972 (.A1(n_6573_o_0),
    .A2(n_6965_o_0),
    .A3(n_6967_o_0),
    .B(n_6971_o_0),
    .Y(n_6972_o_0));
 NOR2xp33_ASAP7_75t_R n_6973 (.A(n_6588_o_0),
    .B(n_6628_o_0),
    .Y(n_6973_o_0));
 OAI211xp5_ASAP7_75t_R n_6974 (.A1(n_6630_o_0),
    .A2(n_6691_o_0),
    .B(n_6624_o_0),
    .C(n_6664_o_0),
    .Y(n_6974_o_0));
 OAI31xp33_ASAP7_75t_R n_6975 (.A1(n_6633_o_0),
    .A2(n_6718_o_0),
    .A3(n_6973_o_0),
    .B(n_6974_o_0),
    .Y(n_6975_o_0));
 NAND2xp33_ASAP7_75t_R n_6976 (.A(n_6831_o_0),
    .B(n_6953_o_0),
    .Y(n_6976_o_0));
 AOI31xp33_ASAP7_75t_R n_6977 (.A1(n_6666_o_0),
    .A2(n_6630_o_0),
    .A3(n_6602_o_0),
    .B(n_6729_o_0),
    .Y(n_6977_o_0));
 AO22x1_ASAP7_75t_R n_6978 (.A1(n_6729_o_0),
    .A2(n_6975_o_0),
    .B1(n_6976_o_0),
    .B2(n_6977_o_0),
    .Y(n_6978_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6979 (.A1(n_6686_o_0),
    .A2(n_6685_o_0),
    .B(n_6624_o_0),
    .C(n_6625_o_0),
    .Y(n_6979_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6980 (.A1(n_6661_o_0),
    .A2(n_6806_o_0),
    .B(n_6777_o_0),
    .C(n_6673_o_0),
    .Y(n_6980_o_0));
 AOI21xp33_ASAP7_75t_R n_6981 (.A1(n_6729_o_0),
    .A2(n_6979_o_0),
    .B(n_6980_o_0),
    .Y(n_6981_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_6982 (.A1(n_6649_o_0),
    .A2(n_6978_o_0),
    .B(n_6679_o_0),
    .C(n_6565_o_0),
    .D(n_6981_o_0),
    .Y(n_6982_o_0));
 AOI211xp5_ASAP7_75t_R n_6983 (.A1(n_6979_o_0),
    .A2(n_6729_o_0),
    .B(n_6980_o_0),
    .C(n_6565_o_0),
    .Y(n_6983_o_0));
 AOI211xp5_ASAP7_75t_R n_6984 (.A1(n_6972_o_0),
    .A2(n_6679_o_0),
    .B(n_6982_o_0),
    .C(n_6983_o_0),
    .Y(n_6984_o_0));
 AOI21xp33_ASAP7_75t_R n_6985 (.A1(n_6962_o_0),
    .A2(n_6708_o_0),
    .B(n_6984_o_0),
    .Y(n_6985_o_0));
 NOR3xp33_ASAP7_75t_R n_6986 (.A(n_6915_o_0),
    .B(n_6899_o_0),
    .C(n_6573_o_0),
    .Y(n_6986_o_0));
 AOI31xp33_ASAP7_75t_R n_6987 (.A1(n_6769_o_0),
    .A2(n_6963_o_0),
    .A3(n_6573_o_0),
    .B(n_6986_o_0),
    .Y(n_6987_o_0));
 AOI211xp5_ASAP7_75t_R n_6988 (.A1(net55),
    .A2(n_6628_o_0),
    .B(n_6666_o_0),
    .C(n_6603_o_0),
    .Y(n_6988_o_0));
 AOI31xp33_ASAP7_75t_R n_6989 (.A1(n_6666_o_0),
    .A2(n_6699_o_0),
    .A3(n_6698_o_0),
    .B(n_6988_o_0),
    .Y(n_6989_o_0));
 AND3x1_ASAP7_75t_R n_6990 (.A(n_6799_o_0),
    .B(n_6670_o_0),
    .C(n_6624_o_0),
    .Y(n_6990_o_0));
 OAI21xp33_ASAP7_75t_R n_6991 (.A1(n_6724_o_0),
    .A2(n_6990_o_0),
    .B(n_6557_o_0),
    .Y(n_6991_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_6992 (.A1(n_6573_o_0),
    .A2(n_6989_o_0),
    .B(n_6991_o_0),
    .C(n_6697_o_0),
    .Y(n_6992_o_0));
 AOI21xp33_ASAP7_75t_R n_6993 (.A1(n_6987_o_0),
    .A2(n_6729_o_0),
    .B(n_6992_o_0),
    .Y(n_6993_o_0));
 AOI32xp33_ASAP7_75t_R n_6994 (.A1(n_6633_o_0),
    .A2(n_6713_o_0),
    .A3(net55),
    .B1(n_6969_o_0),
    .B2(n_6855_o_0),
    .Y(n_6994_o_0));
 NOR2xp33_ASAP7_75t_R n_6995 (.A(n_6630_o_0),
    .B(n_6644_o_0),
    .Y(n_6995_o_0));
 OAI31xp33_ASAP7_75t_R n_6996 (.A1(n_6661_o_0),
    .A2(n_6995_o_0),
    .A3(n_6641_o_0),
    .B(n_6875_o_0),
    .Y(n_6996_o_0));
 AOI22xp33_ASAP7_75t_R n_6997 (.A1(n_6994_o_0),
    .A2(n_6649_o_0),
    .B1(n_6659_o_0),
    .B2(n_6996_o_0),
    .Y(n_6997_o_0));
 AOI21xp33_ASAP7_75t_R n_6998 (.A1(n_6601_o_0),
    .A2(n_6633_o_0),
    .B(n_6957_o_0),
    .Y(n_6998_o_0));
 AOI21xp33_ASAP7_75t_R n_6999 (.A1(n_6624_o_0),
    .A2(n_6757_o_0),
    .B(n_6659_o_0),
    .Y(n_6999_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7000 (.A1(n_6783_o_0),
    .A2(n_6973_o_0),
    .B(n_6999_o_0),
    .C(n_6558_o_0),
    .Y(n_7000_o_0));
 OAI21xp33_ASAP7_75t_R n_7001 (.A1(n_6649_o_0),
    .A2(n_6998_o_0),
    .B(n_7000_o_0),
    .Y(n_7001_o_0));
 OAI21xp33_ASAP7_75t_R n_7002 (.A1(n_6730_o_0),
    .A2(n_6997_o_0),
    .B(n_7001_o_0),
    .Y(n_7002_o_0));
 AO21x1_ASAP7_75t_R n_7003 (.A1(n_7002_o_0),
    .A2(n_6657_o_0),
    .B(n_6707_o_0),
    .Y(n_7003_o_0));
 OAI211xp5_ASAP7_75t_R n_7004 (.A1(n_6601_o_0),
    .A2(net55),
    .B(n_6699_o_0),
    .C(n_6666_o_0),
    .Y(n_7004_o_0));
 OAI21xp33_ASAP7_75t_R n_7005 (.A1(n_6669_o_0),
    .A2(n_6813_o_0),
    .B(n_7004_o_0),
    .Y(n_7005_o_0));
 NAND3xp33_ASAP7_75t_R n_7006 (.A(n_6624_o_0),
    .B(n_6691_o_0),
    .C(net55),
    .Y(n_7006_o_0));
 OAI311xp33_ASAP7_75t_R n_7007 (.A1(n_6633_o_0),
    .A2(n_6784_o_0),
    .A3(n_6662_o_0),
    .B1(n_7006_o_0),
    .C1(n_6558_o_0),
    .Y(n_7007_o_0));
 OAI21xp33_ASAP7_75t_R n_7008 (.A1(n_6729_o_0),
    .A2(n_7005_o_0),
    .B(n_7007_o_0),
    .Y(n_7008_o_0));
 NAND3xp33_ASAP7_75t_R n_7009 (.A(n_6725_o_0),
    .B(n_6671_o_0),
    .C(n_6624_o_0),
    .Y(n_7009_o_0));
 OAI31xp33_ASAP7_75t_R n_7010 (.A1(n_6633_o_0),
    .A2(n_6825_o_0),
    .A3(n_6826_o_0),
    .B(n_7009_o_0),
    .Y(n_7010_o_0));
 AOI21xp33_ASAP7_75t_R n_7011 (.A1(n_6629_o_0),
    .A2(n_6634_o_0),
    .B(n_6729_o_0),
    .Y(n_7011_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7012 (.A1(n_6588_o_0),
    .A2(n_6661_o_0),
    .B(n_7011_o_0),
    .C(n_6573_o_0),
    .Y(n_7012_o_0));
 OAI21xp33_ASAP7_75t_R n_7013 (.A1(n_6557_o_0),
    .A2(n_7010_o_0),
    .B(n_7012_o_0),
    .Y(n_7013_o_0));
 OAI21xp33_ASAP7_75t_R n_7014 (.A1(n_6673_o_0),
    .A2(n_7008_o_0),
    .B(n_7013_o_0),
    .Y(n_7014_o_0));
 OAI21xp33_ASAP7_75t_R n_7015 (.A1(n_6630_o_0),
    .A2(n_6806_o_0),
    .B(n_6633_o_0),
    .Y(n_7015_o_0));
 NAND2xp33_ASAP7_75t_R n_7016 (.A(n_6712_o_0),
    .B(n_7015_o_0),
    .Y(n_7016_o_0));
 AOI31xp33_ASAP7_75t_R n_7017 (.A1(n_6630_o_0),
    .A2(n_6640_o_0),
    .A3(n_6637_o_0),
    .B(n_6633_o_0),
    .Y(n_7017_o_0));
 AOI21xp33_ASAP7_75t_R n_7018 (.A1(n_7017_o_0),
    .A2(n_6799_o_0),
    .B(n_6557_o_0),
    .Y(n_7018_o_0));
 OAI21xp33_ASAP7_75t_R n_7019 (.A1(n_6692_o_0),
    .A2(n_6813_o_0),
    .B(n_7018_o_0),
    .Y(n_7019_o_0));
 OAI211xp5_ASAP7_75t_R n_7020 (.A1(n_6729_o_0),
    .A2(n_7016_o_0),
    .B(n_7019_o_0),
    .C(n_6649_o_0),
    .Y(n_7020_o_0));
 INVx1_ASAP7_75t_R n_7021 (.A(n_6838_o_0),
    .Y(n_7021_o_0));
 AOI21xp33_ASAP7_75t_R n_7022 (.A1(n_6624_o_0),
    .A2(n_7021_o_0),
    .B(n_6729_o_0),
    .Y(n_7022_o_0));
 OAI21xp33_ASAP7_75t_R n_7023 (.A1(n_6784_o_0),
    .A2(n_6719_o_0),
    .B(n_7022_o_0),
    .Y(n_7023_o_0));
 AOI21xp33_ASAP7_75t_R n_7024 (.A1(n_6624_o_0),
    .A2(n_6691_o_0),
    .B(n_6557_o_0),
    .Y(n_7024_o_0));
 OAI21xp33_ASAP7_75t_R n_7025 (.A1(n_6633_o_0),
    .A2(n_6784_o_0),
    .B(n_7024_o_0),
    .Y(n_7025_o_0));
 NAND3xp33_ASAP7_75t_R n_7026 (.A(n_7023_o_0),
    .B(n_7025_o_0),
    .C(n_6659_o_0),
    .Y(n_7026_o_0));
 NAND3xp33_ASAP7_75t_R n_7027 (.A(n_7020_o_0),
    .B(n_7026_o_0),
    .C(n_6674_o_0),
    .Y(n_7027_o_0));
 OAI211xp5_ASAP7_75t_R n_7028 (.A1(n_7014_o_0),
    .A2(n_6657_o_0),
    .B(n_6707_o_0),
    .C(n_7027_o_0),
    .Y(n_7028_o_0));
 OAI21xp33_ASAP7_75t_R n_7029 (.A1(n_6993_o_0),
    .A2(n_7003_o_0),
    .B(n_7028_o_0),
    .Y(n_7029_o_0));
 AOI21xp33_ASAP7_75t_R n_7030 (.A1(n_6588_o_0),
    .A2(net55),
    .B(n_6920_o_0),
    .Y(n_7030_o_0));
 AOI211xp5_ASAP7_75t_R n_7031 (.A1(n_6661_o_0),
    .A2(n_6824_o_0),
    .B(n_7030_o_0),
    .C(n_6673_o_0),
    .Y(n_7031_o_0));
 OAI21xp33_ASAP7_75t_R n_7032 (.A1(n_6756_o_0),
    .A2(n_6624_o_0),
    .B(n_7031_o_0),
    .Y(n_7032_o_0));
 AOI21xp33_ASAP7_75t_R n_7033 (.A1(n_6630_o_0),
    .A2(n_6684_o_0),
    .B(n_6778_o_0),
    .Y(n_7033_o_0));
 AOI21xp33_ASAP7_75t_R n_7034 (.A1(net55),
    .A2(n_6691_o_0),
    .B(n_6949_o_0),
    .Y(n_7034_o_0));
 OAI21xp33_ASAP7_75t_R n_7035 (.A1(n_7033_o_0),
    .A2(n_7034_o_0),
    .B(n_6673_o_0),
    .Y(n_7035_o_0));
 NAND3xp33_ASAP7_75t_R n_7036 (.A(n_7032_o_0),
    .B(n_7035_o_0),
    .C(n_6558_o_0),
    .Y(n_7036_o_0));
 AOI21xp33_ASAP7_75t_R n_7037 (.A1(n_6601_o_0),
    .A2(n_6588_o_0),
    .B(n_6890_o_0),
    .Y(n_7037_o_0));
 AOI31xp33_ASAP7_75t_R n_7038 (.A1(n_6628_o_0),
    .A2(n_6661_o_0),
    .A3(n_6673_o_0),
    .B(n_7037_o_0),
    .Y(n_7038_o_0));
 OAI21xp33_ASAP7_75t_R n_7039 (.A1(n_6633_o_0),
    .A2(n_6773_o_0),
    .B(n_6920_o_0),
    .Y(n_7039_o_0));
 OAI21xp33_ASAP7_75t_R n_7040 (.A1(n_6666_o_0),
    .A2(n_6645_o_0),
    .B(n_7039_o_0),
    .Y(n_7040_o_0));
 AOI21xp33_ASAP7_75t_R n_7041 (.A1(n_6573_o_0),
    .A2(n_7040_o_0),
    .B(n_6558_o_0),
    .Y(n_7041_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7042 (.A1(n_7037_o_0),
    .A2(n_6649_o_0),
    .B(n_7038_o_0),
    .C(n_7041_o_0),
    .Y(n_7042_o_0));
 AOI211xp5_ASAP7_75t_R n_7043 (.A1(n_6713_o_0),
    .A2(net55),
    .B(n_6573_o_0),
    .C(n_6838_o_0),
    .Y(n_7043_o_0));
 AND4x1_ASAP7_75t_R n_7044 (.A(n_6698_o_0),
    .B(n_6615_o_0),
    .C(n_6659_o_0),
    .D(n_6624_o_0),
    .Y(n_7044_o_0));
 AOI21xp33_ASAP7_75t_R n_7045 (.A1(n_6601_o_0),
    .A2(n_6756_o_0),
    .B(n_6666_o_0),
    .Y(n_7045_o_0));
 OA21x2_ASAP7_75t_R n_7046 (.A1(n_6749_o_0),
    .A2(n_7045_o_0),
    .B(n_6649_o_0),
    .Y(n_7046_o_0));
 AOI211xp5_ASAP7_75t_R n_7047 (.A1(n_7043_o_0),
    .A2(n_6666_o_0),
    .B(n_7044_o_0),
    .C(n_7046_o_0),
    .Y(n_7047_o_0));
 OAI21xp33_ASAP7_75t_R n_7048 (.A1(n_6630_o_0),
    .A2(n_6644_o_0),
    .B(n_7017_o_0),
    .Y(n_7048_o_0));
 OAI31xp33_ASAP7_75t_R n_7049 (.A1(n_6661_o_0),
    .A2(n_6669_o_0),
    .A3(n_6718_o_0),
    .B(n_7048_o_0),
    .Y(n_7049_o_0));
 OAI31xp33_ASAP7_75t_R n_7050 (.A1(n_6673_o_0),
    .A2(n_6845_o_0),
    .A3(n_6923_o_0),
    .B(n_6730_o_0),
    .Y(n_7050_o_0));
 AOI21xp33_ASAP7_75t_R n_7051 (.A1(n_6659_o_0),
    .A2(n_7049_o_0),
    .B(n_7050_o_0),
    .Y(n_7051_o_0));
 AOI211xp5_ASAP7_75t_R n_7052 (.A1(n_7047_o_0),
    .A2(n_6558_o_0),
    .B(n_7051_o_0),
    .C(n_6697_o_0),
    .Y(n_7052_o_0));
 AOI31xp33_ASAP7_75t_R n_7053 (.A1(n_6679_o_0),
    .A2(n_7036_o_0),
    .A3(n_7042_o_0),
    .B(n_7052_o_0),
    .Y(n_7053_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7054 (.A1(n_6666_o_0),
    .A2(n_6720_o_0),
    .B(n_6854_o_0),
    .C(n_6615_o_0),
    .Y(n_7054_o_0));
 AOI21xp33_ASAP7_75t_R n_7055 (.A1(n_6603_o_0),
    .A2(n_6633_o_0),
    .B(n_6601_o_0),
    .Y(n_7055_o_0));
 AOI211xp5_ASAP7_75t_R n_7056 (.A1(n_6603_o_0),
    .A2(net55),
    .B(n_7055_o_0),
    .C(n_6649_o_0),
    .Y(n_7056_o_0));
 AOI211xp5_ASAP7_75t_R n_7057 (.A1(n_7054_o_0),
    .A2(n_6573_o_0),
    .B(n_6558_o_0),
    .C(n_7056_o_0),
    .Y(n_7057_o_0));
 OAI21xp33_ASAP7_75t_R n_7058 (.A1(n_6825_o_0),
    .A2(n_6719_o_0),
    .B(n_6573_o_0),
    .Y(n_7058_o_0));
 AOI21xp33_ASAP7_75t_R n_7059 (.A1(n_6624_o_0),
    .A2(n_6762_o_0),
    .B(n_7058_o_0),
    .Y(n_7059_o_0));
 AOI211xp5_ASAP7_75t_R n_7060 (.A1(n_6779_o_0),
    .A2(n_6661_o_0),
    .B(n_6915_o_0),
    .C(n_6573_o_0),
    .Y(n_7060_o_0));
 OAI31xp33_ASAP7_75t_R n_7061 (.A1(n_6557_o_0),
    .A2(n_7059_o_0),
    .A3(n_7060_o_0),
    .B(n_6679_o_0),
    .Y(n_7061_o_0));
 AOI21xp33_ASAP7_75t_R n_7062 (.A1(n_6628_o_0),
    .A2(n_6630_o_0),
    .B(n_6761_o_0),
    .Y(n_7062_o_0));
 OAI21xp33_ASAP7_75t_R n_7063 (.A1(n_6661_o_0),
    .A2(n_7062_o_0),
    .B(n_7004_o_0),
    .Y(n_7063_o_0));
 NOR2xp33_ASAP7_75t_R n_7064 (.A(net55),
    .B(n_6689_o_0),
    .Y(n_7064_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7065 (.A1(n_7064_o_0),
    .A2(n_7015_o_0),
    .B(n_6775_o_0),
    .C(n_6659_o_0),
    .Y(n_7065_o_0));
 AOI211xp5_ASAP7_75t_R n_7066 (.A1(n_6673_o_0),
    .A2(n_7063_o_0),
    .B(n_7065_o_0),
    .C(n_6558_o_0),
    .Y(n_7066_o_0));
 INVx1_ASAP7_75t_R n_7067 (.A(n_6703_o_0),
    .Y(n_7067_o_0));
 AOI21xp33_ASAP7_75t_R n_7068 (.A1(n_7067_o_0),
    .A2(n_6976_o_0),
    .B(n_6659_o_0),
    .Y(n_7068_o_0));
 AOI211xp5_ASAP7_75t_R n_7069 (.A1(n_6659_o_0),
    .A2(n_6827_o_0),
    .B(n_7068_o_0),
    .C(n_6730_o_0),
    .Y(n_7069_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7070 (.A1(n_7066_o_0),
    .A2(n_7069_o_0),
    .B(n_6657_o_0),
    .C(n_6708_o_0),
    .Y(n_7070_o_0));
 OAI21xp33_ASAP7_75t_R n_7071 (.A1(n_7057_o_0),
    .A2(n_7061_o_0),
    .B(n_7070_o_0),
    .Y(n_7071_o_0));
 OAI21xp33_ASAP7_75t_R n_7072 (.A1(n_6565_o_0),
    .A2(n_7053_o_0),
    .B(n_7071_o_0),
    .Y(n_7072_o_0));
 NOR2xp33_ASAP7_75t_R n_7073 (.A(n_6973_o_0),
    .B(n_6823_o_0),
    .Y(n_7073_o_0));
 AOI31xp33_ASAP7_75t_R n_7074 (.A1(n_6624_o_0),
    .A2(n_6699_o_0),
    .A3(n_7021_o_0),
    .B(n_7073_o_0),
    .Y(n_7074_o_0));
 OAI21xp33_ASAP7_75t_R n_7075 (.A1(n_6588_o_0),
    .A2(n_6628_o_0),
    .B(n_6614_o_0),
    .Y(n_7075_o_0));
 NAND3xp33_ASAP7_75t_R n_7076 (.A(n_6909_o_0),
    .B(n_7075_o_0),
    .C(n_6661_o_0),
    .Y(n_7076_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7077 (.A1(n_6691_o_0),
    .A2(net55),
    .B(n_6714_o_0),
    .C(n_7076_o_0),
    .Y(n_7077_o_0));
 OAI22xp33_ASAP7_75t_R n_7078 (.A1(n_7074_o_0),
    .A2(n_6673_o_0),
    .B1(n_7077_o_0),
    .B2(n_6573_o_0),
    .Y(n_7078_o_0));
 NOR3xp33_ASAP7_75t_R n_7079 (.A(n_6624_o_0),
    .B(n_6628_o_0),
    .C(n_6603_o_0),
    .Y(n_7079_o_0));
 OAI211xp5_ASAP7_75t_R n_7080 (.A1(n_6666_o_0),
    .A2(n_6958_o_0),
    .B(n_6774_o_0),
    .C(n_6733_o_0),
    .Y(n_7080_o_0));
 OAI31xp33_ASAP7_75t_R n_7081 (.A1(n_6673_o_0),
    .A2(n_7037_o_0),
    .A3(n_7079_o_0),
    .B(n_7080_o_0),
    .Y(n_7081_o_0));
 OAI21xp33_ASAP7_75t_R n_7082 (.A1(n_6557_o_0),
    .A2(n_7081_o_0),
    .B(n_6679_o_0),
    .Y(n_7082_o_0));
 AOI21xp33_ASAP7_75t_R n_7083 (.A1(n_6557_o_0),
    .A2(n_7078_o_0),
    .B(n_7082_o_0),
    .Y(n_7083_o_0));
 OA21x2_ASAP7_75t_R n_7084 (.A1(n_6718_o_0),
    .A2(n_6783_o_0),
    .B(n_6874_o_0),
    .Y(n_7084_o_0));
 AOI31xp33_ASAP7_75t_R n_7085 (.A1(n_6666_o_0),
    .A2(n_6851_o_0),
    .A3(n_6646_o_0),
    .B(n_6649_o_0),
    .Y(n_7085_o_0));
 OAI21xp33_ASAP7_75t_R n_7086 (.A1(n_6661_o_0),
    .A2(n_6759_o_0),
    .B(n_7085_o_0),
    .Y(n_7086_o_0));
 OAI21xp33_ASAP7_75t_R n_7087 (.A1(n_6673_o_0),
    .A2(n_7084_o_0),
    .B(n_7086_o_0),
    .Y(n_7087_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7088 (.A1(n_6628_o_0),
    .A2(n_6603_o_0),
    .B(n_6630_o_0),
    .C(n_6890_o_0),
    .Y(n_7088_o_0));
 AOI21xp33_ASAP7_75t_R n_7089 (.A1(n_6601_o_0),
    .A2(n_6756_o_0),
    .B(n_6624_o_0),
    .Y(n_7089_o_0));
 OAI21xp33_ASAP7_75t_R n_7090 (.A1(n_6661_o_0),
    .A2(n_6806_o_0),
    .B(n_6733_o_0),
    .Y(n_7090_o_0));
 OAI31xp33_ASAP7_75t_R n_7091 (.A1(n_6673_o_0),
    .A2(n_7088_o_0),
    .A3(n_7089_o_0),
    .B(n_7090_o_0),
    .Y(n_7091_o_0));
 OAI21xp33_ASAP7_75t_R n_7092 (.A1(n_6729_o_0),
    .A2(n_7091_o_0),
    .B(n_6657_o_0),
    .Y(n_7092_o_0));
 AOI21xp33_ASAP7_75t_R n_7093 (.A1(n_6729_o_0),
    .A2(n_7087_o_0),
    .B(n_7092_o_0),
    .Y(n_7093_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7094 (.A1(n_6630_o_0),
    .A2(n_6603_o_0),
    .B(n_6899_o_0),
    .C(n_6807_o_0),
    .Y(n_7094_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7095 (.A1(n_6909_o_0),
    .A2(n_7075_o_0),
    .B(n_6661_o_0),
    .C(n_6730_o_0),
    .Y(n_7095_o_0));
 AOI31xp33_ASAP7_75t_R n_7096 (.A1(n_6666_o_0),
    .A2(n_6671_o_0),
    .A3(n_6698_o_0),
    .B(n_7095_o_0),
    .Y(n_7096_o_0));
 AOI211xp5_ASAP7_75t_R n_7097 (.A1(n_7094_o_0),
    .A2(n_6558_o_0),
    .B(n_6673_o_0),
    .C(n_7096_o_0),
    .Y(n_7097_o_0));
 OAI21xp33_ASAP7_75t_R n_7098 (.A1(net55),
    .A2(n_6806_o_0),
    .B(n_6661_o_0),
    .Y(n_7098_o_0));
 AO21x1_ASAP7_75t_R n_7099 (.A1(n_6976_o_0),
    .A2(n_7098_o_0),
    .B(n_6729_o_0),
    .Y(n_7099_o_0));
 OAI21xp33_ASAP7_75t_R n_7100 (.A1(n_7034_o_0),
    .A2(n_6868_o_0),
    .B(n_6558_o_0),
    .Y(n_7100_o_0));
 AOI21xp33_ASAP7_75t_R n_7101 (.A1(n_7099_o_0),
    .A2(n_7100_o_0),
    .B(n_6649_o_0),
    .Y(n_7101_o_0));
 NOR3xp33_ASAP7_75t_R n_7102 (.A(n_6779_o_0),
    .B(n_6636_o_0),
    .C(n_6633_o_0),
    .Y(n_7102_o_0));
 OAI21xp33_ASAP7_75t_R n_7103 (.A1(n_6761_o_0),
    .A2(n_6693_o_0),
    .B(n_6730_o_0),
    .Y(n_7103_o_0));
 AOI21xp33_ASAP7_75t_R n_7104 (.A1(n_6588_o_0),
    .A2(n_6666_o_0),
    .B(n_7103_o_0),
    .Y(n_7104_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7105 (.A1(n_6624_o_0),
    .A2(n_6698_o_0),
    .B(n_7102_o_0),
    .C(n_6729_o_0),
    .D(n_7104_o_0),
    .Y(n_7105_o_0));
 NAND2xp33_ASAP7_75t_R n_7106 (.A(n_6854_o_0),
    .B(n_6855_o_0),
    .Y(n_7106_o_0));
 OAI31xp33_ASAP7_75t_R n_7107 (.A1(n_6633_o_0),
    .A2(n_6636_o_0),
    .A3(n_6718_o_0),
    .B(n_7106_o_0),
    .Y(n_7107_o_0));
 NAND2xp33_ASAP7_75t_R n_7108 (.A(n_6557_o_0),
    .B(n_7107_o_0),
    .Y(n_7108_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7109 (.A1(n_6666_o_0),
    .A2(n_6689_o_0),
    .B(n_6766_o_0),
    .C(n_6630_o_0),
    .Y(n_7109_o_0));
 OA21x2_ASAP7_75t_R n_7110 (.A1(n_7109_o_0),
    .A2(n_6730_o_0),
    .B(n_6673_o_0),
    .Y(n_7110_o_0));
 AOI22xp33_ASAP7_75t_R n_7111 (.A1(n_7105_o_0),
    .A2(n_6573_o_0),
    .B1(n_7108_o_0),
    .B2(n_7110_o_0),
    .Y(n_7111_o_0));
 OAI321xp33_ASAP7_75t_R n_7112 (.A1(n_6657_o_0),
    .A2(n_7097_o_0),
    .A3(n_7101_o_0),
    .B1(n_7111_o_0),
    .B2(n_6679_o_0),
    .C(n_6707_o_0),
    .Y(n_7112_o_0));
 OAI31xp33_ASAP7_75t_R n_7113 (.A1(n_6565_o_0),
    .A2(n_7083_o_0),
    .A3(n_7093_o_0),
    .B(n_7112_o_0),
    .Y(n_7113_o_0));
 XNOR2xp5_ASAP7_75t_R n_7114 (.A(_01073_),
    .B(_01074_),
    .Y(n_7114_o_0));
 XNOR2xp5_ASAP7_75t_R n_7115 (.A(_01113_),
    .B(n_7114_o_0),
    .Y(n_7115_o_0));
 XOR2xp5_ASAP7_75t_R n_7116 (.A(_01026_),
    .B(_01033_),
    .Y(n_7116_o_0));
 NOR2xp33_ASAP7_75t_R n_7117 (.A(n_7116_o_0),
    .B(n_7115_o_0),
    .Y(n_7117_o_0));
 NOR2xp33_ASAP7_75t_R n_7118 (.A(_00715_),
    .B(net),
    .Y(n_7118_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7119 (.A1(n_7115_o_0),
    .A2(n_7116_o_0),
    .B(n_7117_o_0),
    .C(net),
    .D(n_7118_o_0),
    .Y(n_7119_o_0));
 NOR2xp33_ASAP7_75t_R n_7120 (.A(_00978_),
    .B(n_7119_o_0),
    .Y(n_7120_o_0));
 XOR2xp5_ASAP7_75t_R n_7121 (.A(_01027_),
    .B(_01034_),
    .Y(n_7121_o_0));
 XNOR2xp5_ASAP7_75t_R n_7122 (.A(_01074_),
    .B(_01075_),
    .Y(n_7122_o_0));
 XNOR2xp5_ASAP7_75t_R n_7123 (.A(_01114_),
    .B(n_7122_o_0),
    .Y(n_7123_o_0));
 XNOR2xp5_ASAP7_75t_R n_7124 (.A(n_7121_o_0),
    .B(n_7123_o_0),
    .Y(n_7124_o_0));
 NOR2xp33_ASAP7_75t_R n_7125 (.A(_00714_),
    .B(net),
    .Y(n_7125_o_0));
 AOI21xp33_ASAP7_75t_R n_7126 (.A1(net),
    .A2(n_7124_o_0),
    .B(n_7125_o_0),
    .Y(n_7126_o_0));
 HAxp5_ASAP7_75t_R n_7127 (.A(n_964_o_0),
    .B(n_7126_o_0),
    .CON(n_7127_o_0),
    .SN(n_7127_o_1));
 XNOR2xp5_ASAP7_75t_R n_7128 (.A(_01025_),
    .B(_01032_),
    .Y(n_7128_o_0));
 XNOR2xp5_ASAP7_75t_R n_7129 (.A(_01072_),
    .B(n_7128_o_0),
    .Y(n_7129_o_0));
 XOR2xp5_ASAP7_75t_R n_7130 (.A(n_4804_o_0),
    .B(n_7129_o_0),
    .Y(n_7130_o_0));
 NOR2xp33_ASAP7_75t_R n_7131 (.A(_00716_),
    .B(net),
    .Y(n_7131_o_0));
 AOI21xp33_ASAP7_75t_R n_7132 (.A1(net),
    .A2(n_7130_o_0),
    .B(n_7131_o_0),
    .Y(n_7132_o_0));
 NAND2xp33_ASAP7_75t_R n_7133 (.A(_00977_),
    .B(n_7132_o_0),
    .Y(n_7133_o_0));
 OAI21xp33_ASAP7_75t_R n_7134 (.A1(_00977_),
    .A2(n_7132_o_0),
    .B(n_7133_o_0),
    .Y(n_7134_o_0));
 NOR2xp33_ASAP7_75t_R n_7135 (.A(_00718_),
    .B(_00858_),
    .Y(n_7135_o_0));
 NAND2xp33_ASAP7_75t_R n_7136 (.A(n_3021_o_0),
    .B(n_7135_o_0),
    .Y(n_7136_o_0));
 XNOR2xp5_ASAP7_75t_R n_7137 (.A(_01070_),
    .B(_01075_),
    .Y(n_7137_o_0));
 XNOR2xp5_ASAP7_75t_R n_7138 (.A(n_4837_o_0),
    .B(n_7137_o_0),
    .Y(n_7138_o_0));
 INVx1_ASAP7_75t_R n_7139 (.A(_01023_),
    .Y(n_7139_o_0));
 XNOR2xp5_ASAP7_75t_R n_7140 (.A(n_7139_o_0),
    .B(n_4836_o_0),
    .Y(n_7140_o_0));
 NAND2xp33_ASAP7_75t_R n_7141 (.A(n_7139_o_0),
    .B(n_4844_o_0),
    .Y(n_7141_o_0));
 NAND2xp33_ASAP7_75t_R n_7142 (.A(_01023_),
    .B(n_4836_o_0),
    .Y(n_7142_o_0));
 XOR2xp5_ASAP7_75t_R n_7143 (.A(_01070_),
    .B(_01075_),
    .Y(n_7143_o_0));
 NAND2xp33_ASAP7_75t_R n_7144 (.A(n_4837_o_0),
    .B(n_7143_o_0),
    .Y(n_7144_o_0));
 NAND2xp33_ASAP7_75t_R n_7145 (.A(n_7137_o_0),
    .B(n_4842_o_0),
    .Y(n_7145_o_0));
 AOI22xp33_ASAP7_75t_R n_7146 (.A1(n_7141_o_0),
    .A2(n_7142_o_0),
    .B1(n_7144_o_0),
    .B2(n_7145_o_0),
    .Y(n_7146_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7147 (.A1(n_7138_o_0),
    .A2(n_7140_o_0),
    .B(n_7146_o_0),
    .C(net39),
    .Y(n_7147_o_0));
 NAND2xp33_ASAP7_75t_R n_7148 (.A(n_7136_o_0),
    .B(n_7147_o_0),
    .Y(n_7148_o_0));
 AOI21xp33_ASAP7_75t_R n_7149 (.A1(n_7136_o_0),
    .A2(n_7147_o_0),
    .B(n_874_o_0),
    .Y(n_7149_o_0));
 INVx1_ASAP7_75t_R n_7150 (.A(n_7149_o_0),
    .Y(n_7150_o_0));
 OAI21xp33_ASAP7_75t_R n_7151 (.A1(_00975_),
    .A2(n_7148_o_0),
    .B(n_7150_o_0),
    .Y(n_7151_o_0));
 XNOR2xp5_ASAP7_75t_R n_7152 (.A(_01068_),
    .B(_01075_),
    .Y(n_7152_o_0));
 XOR2xp5_ASAP7_75t_R n_7153 (.A(_01069_),
    .B(_01108_),
    .Y(n_7153_o_0));
 XNOR2xp5_ASAP7_75t_R n_7154 (.A(n_7152_o_0),
    .B(n_7153_o_0),
    .Y(n_7154_o_0));
 XNOR2xp5_ASAP7_75t_R n_7155 (.A(_01021_),
    .B(n_4906_o_0),
    .Y(n_7155_o_0));
 XOR2xp5_ASAP7_75t_R n_7156 (.A(_01068_),
    .B(_01075_),
    .Y(n_7156_o_0));
 NAND2xp33_ASAP7_75t_R n_7157 (.A(n_7156_o_0),
    .B(n_7153_o_0),
    .Y(n_7157_o_0));
 XNOR2xp5_ASAP7_75t_R n_7158 (.A(_01069_),
    .B(_01108_),
    .Y(n_7158_o_0));
 NAND2xp33_ASAP7_75t_R n_7159 (.A(n_7152_o_0),
    .B(n_7158_o_0),
    .Y(n_7159_o_0));
 NAND2xp33_ASAP7_75t_R n_7160 (.A(_01021_),
    .B(n_4928_o_0),
    .Y(n_7160_o_0));
 INVx1_ASAP7_75t_R n_7161 (.A(_01021_),
    .Y(n_7161_o_0));
 NAND2xp33_ASAP7_75t_R n_7162 (.A(n_7161_o_0),
    .B(n_4906_o_0),
    .Y(n_7162_o_0));
 AOI22xp33_ASAP7_75t_R n_7163 (.A1(n_7157_o_0),
    .A2(n_7159_o_0),
    .B1(n_7160_o_0),
    .B2(n_7162_o_0),
    .Y(n_7163_o_0));
 NOR2xp33_ASAP7_75t_R n_7164 (.A(_00559_),
    .B(_00858_),
    .Y(n_7164_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7165 (.A1(n_7154_o_0),
    .A2(n_7155_o_0),
    .B(n_7163_o_0),
    .C(_00858_),
    .D(n_7164_o_0),
    .Y(n_7165_o_0));
 NAND2xp33_ASAP7_75t_R n_7166 (.A(_00973_),
    .B(n_7165_o_0),
    .Y(n_7166_o_0));
 NAND2xp33_ASAP7_75t_R n_7167 (.A(_01035_),
    .B(_01107_),
    .Y(n_7167_o_0));
 OA21x2_ASAP7_75t_R n_7168 (.A1(_01035_),
    .A2(_01107_),
    .B(n_7167_o_0),
    .Y(n_7168_o_0));
 OAI211xp5_ASAP7_75t_R n_7169 (.A1(_01035_),
    .A2(_01107_),
    .B(n_7167_o_0),
    .C(n_4922_o_0),
    .Y(n_7169_o_0));
 OAI21xp33_ASAP7_75t_R n_7170 (.A1(n_4922_o_0),
    .A2(n_7168_o_0),
    .B(n_7169_o_0),
    .Y(n_7170_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7171 (.A1(_01035_),
    .A2(_01107_),
    .B(n_7167_o_0),
    .C(n_4922_o_0),
    .Y(n_7171_o_0));
 AOI211xp5_ASAP7_75t_R n_7172 (.A1(n_7168_o_0),
    .A2(n_4922_o_0),
    .B(n_7156_o_0),
    .C(n_7171_o_0),
    .Y(n_7172_o_0));
 NOR2xp33_ASAP7_75t_R n_7173 (.A(_00560_),
    .B(_00858_),
    .Y(n_7173_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7174 (.A1(n_7156_o_0),
    .A2(n_7170_o_0),
    .B(n_7172_o_0),
    .C(net39),
    .D(n_7173_o_0),
    .Y(n_7174_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7175 (.A1(n_7168_o_0),
    .A2(n_4922_o_0),
    .B(n_7171_o_0),
    .C(n_7156_o_0),
    .Y(n_7175_o_0));
 OAI211xp5_ASAP7_75t_R n_7176 (.A1(n_7168_o_0),
    .A2(n_4922_o_0),
    .B(n_7169_o_0),
    .C(n_7152_o_0),
    .Y(n_7176_o_0));
 INVx1_ASAP7_75t_R n_7177 (.A(n_7173_o_0),
    .Y(n_7177_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7178 (.A1(n_7175_o_0),
    .A2(n_7176_o_0),
    .B(net1),
    .C(n_7177_o_0),
    .D(_00972_),
    .Y(n_7178_o_0));
 AOI21x1_ASAP7_75t_R n_7179 (.A1(_00972_),
    .A2(n_7174_o_0),
    .B(n_7178_o_0),
    .Y(n_7179_o_0));
 OAI211xp5_ASAP7_75t_R n_7180 (.A1(_00973_),
    .A2(n_7165_o_0),
    .B(n_7166_o_0),
    .C(n_7179_o_0),
    .Y(n_7180_o_0));
 NOR2xp33_ASAP7_75t_R n_7181 (.A(_00973_),
    .B(n_7165_o_0),
    .Y(n_7181_o_0));
 AO21x1_ASAP7_75t_R n_7182 (.A1(_00972_),
    .A2(n_7174_o_0),
    .B(n_7178_o_0),
    .Y(n_7182_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7183 (.A1(_00973_),
    .A2(n_7165_o_0),
    .B(n_7181_o_0),
    .C(n_7182_o_0),
    .Y(n_7183_o_0));
 INVx1_ASAP7_75t_R n_7184 (.A(_01022_),
    .Y(n_7184_o_0));
 NAND2xp33_ASAP7_75t_R n_7185 (.A(n_7184_o_0),
    .B(n_4863_o_0),
    .Y(n_7185_o_0));
 INVx1_ASAP7_75t_R n_7186 (.A(n_7185_o_0),
    .Y(n_7186_o_0));
 NOR2xp33_ASAP7_75t_R n_7187 (.A(n_7184_o_0),
    .B(n_4863_o_0),
    .Y(n_7187_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7188 (.A1(n_4863_o_0),
    .A2(n_7184_o_0),
    .B(n_7187_o_0),
    .C(n_4926_o_0),
    .Y(n_7188_o_0));
 OAI31xp33_ASAP7_75t_R n_7189 (.A1(n_7186_o_0),
    .A2(n_7187_o_0),
    .A3(n_4926_o_0),
    .B(n_7188_o_0),
    .Y(n_7189_o_0));
 NOR2xp33_ASAP7_75t_R n_7190 (.A(_00562_),
    .B(_00858_),
    .Y(n_7190_o_0));
 AOI21xp33_ASAP7_75t_R n_7191 (.A1(_00858_),
    .A2(n_7189_o_0),
    .B(n_7190_o_0),
    .Y(n_7191_o_0));
 INVx1_ASAP7_75t_R n_7192 (.A(_00974_),
    .Y(n_7192_o_0));
 OAI211xp5_ASAP7_75t_R n_7193 (.A1(n_4863_o_0),
    .A2(n_7184_o_0),
    .B(n_7185_o_0),
    .C(n_4912_o_0),
    .Y(n_7193_o_0));
 INVx1_ASAP7_75t_R n_7194 (.A(n_7190_o_0),
    .Y(n_7194_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7195 (.A1(n_7193_o_0),
    .A2(n_7188_o_0),
    .B(n_3021_o_0),
    .C(n_7194_o_0),
    .D(n_7192_o_0),
    .Y(n_7195_o_0));
 AO21x2_ASAP7_75t_R n_7196 (.A1(n_7191_o_0),
    .A2(n_7192_o_0),
    .B(n_7195_o_0),
    .Y(n_7196_o_0));
 AOI21xp33_ASAP7_75t_R n_7197 (.A1(n_7180_o_0),
    .A2(n_7183_o_0),
    .B(n_7196_o_0),
    .Y(n_7197_o_0));
 INVx1_ASAP7_75t_R n_7198 (.A(n_7197_o_0),
    .Y(n_7198_o_0));
 AOI21x1_ASAP7_75t_R n_7199 (.A1(_00973_),
    .A2(n_7165_o_0),
    .B(n_7181_o_0),
    .Y(n_7199_o_0));
 AOI21x1_ASAP7_75t_R n_7200 (.A1(n_7192_o_0),
    .A2(n_7191_o_0),
    .B(n_7195_o_0),
    .Y(n_7200_o_0));
 OAI21x1_ASAP7_75t_R n_7201 (.A1(_00973_),
    .A2(n_7165_o_0),
    .B(n_7166_o_0),
    .Y(n_7201_o_0));
 OAI21x1_ASAP7_75t_R n_7202 (.A1(n_7182_o_0),
    .A2(n_7201_o_0),
    .B(n_7183_o_0),
    .Y(n_7202_o_0));
 AO21x1_ASAP7_75t_R n_7203 (.A1(n_7138_o_0),
    .A2(n_7140_o_0),
    .B(n_7146_o_0),
    .Y(n_7203_o_0));
 AOI211xp5_ASAP7_75t_R n_7204 (.A1(n_7203_o_0),
    .A2(net39),
    .B(n_874_o_0),
    .C(n_7135_o_0),
    .Y(n_7204_o_0));
 AO21x1_ASAP7_75t_R n_7205 (.A1(n_874_o_0),
    .A2(n_7148_o_0),
    .B(n_7204_o_0),
    .Y(n_7205_o_0));
 OAI21xp33_ASAP7_75t_R n_7206 (.A1(n_7200_o_0),
    .A2(n_7202_o_0),
    .B(n_7205_o_0),
    .Y(n_7206_o_0));
 XNOR2xp5_ASAP7_75t_R n_7207 (.A(_01024_),
    .B(n_4958_o_0),
    .Y(n_7207_o_0));
 XNOR2xp5_ASAP7_75t_R n_7208 (.A(_01071_),
    .B(_01075_),
    .Y(n_7208_o_0));
 XNOR2xp5_ASAP7_75t_R n_7209 (.A(n_4959_o_0),
    .B(n_7208_o_0),
    .Y(n_7209_o_0));
 XOR2xp5_ASAP7_75t_R n_7210 (.A(n_7207_o_0),
    .B(n_7209_o_0),
    .Y(n_7210_o_0));
 NOR2xp33_ASAP7_75t_R n_7211 (.A(_00717_),
    .B(_00858_),
    .Y(n_7211_o_0));
 AOI21xp33_ASAP7_75t_R n_7212 (.A1(net39),
    .A2(n_7210_o_0),
    .B(n_7211_o_0),
    .Y(n_7212_o_0));
 XNOR2xp5_ASAP7_75t_R n_7213 (.A(n_825_o_0),
    .B(n_7212_o_0),
    .Y(n_7213_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7214 (.A1(net79),
    .A2(net46),
    .B(n_7206_o_0),
    .C(n_7213_o_0),
    .Y(n_7214_o_0));
 AO21x1_ASAP7_75t_R n_7215 (.A1(n_7151_o_0),
    .A2(n_7198_o_0),
    .B(n_7214_o_0),
    .Y(n_7215_o_0));
 NAND2x1_ASAP7_75t_R n_7216 (.A(n_7182_o_0),
    .B(n_7201_o_0),
    .Y(n_7216_o_0));
 NAND3xp33_ASAP7_75t_R n_7217 (.A(n_7216_o_0),
    .B(n_7196_o_0),
    .C(n_7205_o_0),
    .Y(n_7217_o_0));
 INVx1_ASAP7_75t_R n_7218 (.A(n_7217_o_0),
    .Y(n_7218_o_0));
 AOI21x1_ASAP7_75t_R n_7219 (.A1(n_874_o_0),
    .A2(n_7148_o_0),
    .B(n_7204_o_0),
    .Y(n_7219_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7220 (.A1(_00973_),
    .A2(n_7165_o_0),
    .B(n_7181_o_0),
    .C(n_7179_o_0),
    .Y(n_7220_o_0));
 INVx1_ASAP7_75t_R n_7221 (.A(n_7220_o_0),
    .Y(n_7221_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7222 (.A1(_00973_),
    .A2(n_7165_o_0),
    .B(n_7166_o_0),
    .C(n_7179_o_0),
    .Y(n_7222_o_0));
 AOI211xp5_ASAP7_75t_R n_7223 (.A1(_00973_),
    .A2(n_7165_o_0),
    .B(n_7181_o_0),
    .C(n_7182_o_0),
    .Y(n_7223_o_0));
 AOI31xp67_ASAP7_75t_R n_7224 (.A1(n_874_o_0),
    .A2(n_7136_o_0),
    .A3(n_7147_o_0),
    .B(n_7149_o_0),
    .Y(n_7224_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7225 (.A1(n_7222_o_0),
    .A2(n_7223_o_0),
    .B(n_7196_o_0),
    .C(n_7224_o_0),
    .Y(n_7225_o_0));
 OAI21xp33_ASAP7_75t_R n_7226 (.A1(n_7216_o_0),
    .A2(n_7196_o_0),
    .B(n_7225_o_0),
    .Y(n_7226_o_0));
 OAI31xp33_ASAP7_75t_R n_7227 (.A1(n_7219_o_0),
    .A2(n_7221_o_0),
    .A3(n_7196_o_0),
    .B(n_7226_o_0),
    .Y(n_7227_o_0));
 NAND2xp33_ASAP7_75t_R n_7228 (.A(_00976_),
    .B(n_7212_o_0),
    .Y(n_7228_o_0));
 OAI21xp33_ASAP7_75t_R n_7229 (.A1(_00976_),
    .A2(n_7212_o_0),
    .B(n_7228_o_0),
    .Y(n_7229_o_0));
 OAI21xp33_ASAP7_75t_R n_7230 (.A1(n_7218_o_0),
    .A2(n_7227_o_0),
    .B(n_7229_o_0),
    .Y(n_7230_o_0));
 NOR2xp33_ASAP7_75t_R n_7231 (.A(n_7179_o_0),
    .B(n_7201_o_0),
    .Y(n_7231_o_0));
 NOR2xp33_ASAP7_75t_R n_7232 (.A(n_7182_o_0),
    .B(n_7196_o_0),
    .Y(n_7232_o_0));
 NAND2xp33_ASAP7_75t_R n_7233 (.A(n_7179_o_0),
    .B(n_7196_o_0),
    .Y(n_7233_o_0));
 NAND2xp33_ASAP7_75t_R n_7234 (.A(n_7182_o_0),
    .B(n_7201_o_0),
    .Y(n_7234_o_0));
 NAND3xp33_ASAP7_75t_R n_7235 (.A(n_7233_o_0),
    .B(n_7234_o_0),
    .C(n_7205_o_0),
    .Y(n_7235_o_0));
 OAI31xp33_ASAP7_75t_R n_7236 (.A1(n_7224_o_0),
    .A2(n_7231_o_0),
    .A3(n_7232_o_0),
    .B(n_7235_o_0),
    .Y(n_7236_o_0));
 XNOR2xp5_ASAP7_75t_R n_7237 (.A(n_7207_o_0),
    .B(n_7209_o_0),
    .Y(n_7237_o_0));
 INVx1_ASAP7_75t_R n_7238 (.A(n_7211_o_0),
    .Y(n_7238_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7239 (.A1(net1),
    .A2(n_7237_o_0),
    .B(n_7238_o_0),
    .C(n_825_o_0),
    .Y(n_7239_o_0));
 AOI21xp5_ASAP7_75t_R n_7240 (.A1(n_825_o_0),
    .A2(n_7212_o_0),
    .B(n_7239_o_0),
    .Y(n_7240_o_0));
 INVx2_ASAP7_75t_R n_7241 (.A(n_7240_o_0),
    .Y(n_7241_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7242 (.A1(n_7183_o_0),
    .A2(n_7180_o_0),
    .B(n_7200_o_0),
    .C(n_7224_o_0),
    .Y(n_7242_o_0));
 NOR3xp33_ASAP7_75t_R n_7243 (.A(n_7196_o_0),
    .B(n_7201_o_0),
    .C(n_7182_o_0),
    .Y(n_7243_o_0));
 AOI21xp33_ASAP7_75t_R n_7244 (.A1(n_7179_o_0),
    .A2(n_7201_o_0),
    .B(n_7200_o_0),
    .Y(n_7244_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7245 (.A1(n_7216_o_0),
    .A2(net46),
    .B(n_7244_o_0),
    .C(n_7219_o_0),
    .Y(n_7245_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7246 (.A1(n_7242_o_0),
    .A2(n_7243_o_0),
    .B(n_7245_o_0),
    .C(n_7241_o_0),
    .Y(n_7246_o_0));
 AOI211xp5_ASAP7_75t_R n_7247 (.A1(n_7236_o_0),
    .A2(n_7241_o_0),
    .B(n_7134_o_0),
    .C(n_7246_o_0),
    .Y(n_7247_o_0));
 AOI31xp33_ASAP7_75t_R n_7248 (.A1(n_7134_o_0),
    .A2(n_7215_o_0),
    .A3(n_7230_o_0),
    .B(n_7247_o_0),
    .Y(n_7248_o_0));
 AOI21xp33_ASAP7_75t_R n_7249 (.A1(n_7200_o_0),
    .A2(n_7220_o_0),
    .B(n_7224_o_0),
    .Y(n_7249_o_0));
 NOR2xp33_ASAP7_75t_R n_7250 (.A(n_7200_o_0),
    .B(n_7179_o_0),
    .Y(n_7250_o_0));
 NAND2xp33_ASAP7_75t_R n_7251 (.A(n_7199_o_0),
    .B(n_7250_o_0),
    .Y(n_7251_o_0));
 AOI21xp33_ASAP7_75t_R n_7252 (.A1(n_7249_o_0),
    .A2(n_7251_o_0),
    .B(n_7241_o_0),
    .Y(n_7252_o_0));
 OAI31xp33_ASAP7_75t_R n_7253 (.A1(n_7216_o_0),
    .A2(net46),
    .A3(n_7219_o_0),
    .B(n_7252_o_0),
    .Y(n_7253_o_0));
 OAI21xp33_ASAP7_75t_R n_7254 (.A1(n_7196_o_0),
    .A2(n_7220_o_0),
    .B(n_7205_o_0),
    .Y(n_7254_o_0));
 INVx1_ASAP7_75t_R n_7255 (.A(n_7254_o_0),
    .Y(n_7255_o_0));
 AOI21xp33_ASAP7_75t_R n_7256 (.A1(n_7251_o_0),
    .A2(n_7255_o_0),
    .B(n_7229_o_0),
    .Y(n_7256_o_0));
 OAI31xp33_ASAP7_75t_R n_7257 (.A1(n_7216_o_0),
    .A2(net46),
    .A3(n_7224_o_0),
    .B(n_7256_o_0),
    .Y(n_7257_o_0));
 NAND2xp33_ASAP7_75t_R n_7258 (.A(n_7253_o_0),
    .B(n_7257_o_0),
    .Y(n_7258_o_0));
 NAND2xp33_ASAP7_75t_R n_7259 (.A(n_900_o_0),
    .B(n_7132_o_0),
    .Y(n_7259_o_0));
 OAI21xp33_ASAP7_75t_R n_7260 (.A1(n_7132_o_0),
    .A2(n_900_o_0),
    .B(n_7259_o_0),
    .Y(n_7260_o_0));
 INVx1_ASAP7_75t_R n_7261 (.A(n_7260_o_0),
    .Y(n_7261_o_0));
 NOR2xp33_ASAP7_75t_R n_7262 (.A(n_7179_o_0),
    .B(n_7201_o_0),
    .Y(n_7262_o_0));
 NOR2xp33_ASAP7_75t_R n_7263 (.A(n_7200_o_0),
    .B(n_7201_o_0),
    .Y(n_7263_o_0));
 AOI21xp33_ASAP7_75t_R n_7264 (.A1(n_7182_o_0),
    .A2(n_7263_o_0),
    .B(n_7151_o_0),
    .Y(n_7264_o_0));
 OAI21xp33_ASAP7_75t_R n_7265 (.A1(n_7196_o_0),
    .A2(n_7262_o_0),
    .B(n_7264_o_0),
    .Y(n_7265_o_0));
 NOR2xp33_ASAP7_75t_R n_7266 (.A(n_7179_o_0),
    .B(n_7199_o_0),
    .Y(n_7266_o_0));
 NOR2xp33_ASAP7_75t_R n_7267 (.A(n_7196_o_0),
    .B(n_7151_o_0),
    .Y(n_7267_o_0));
 NAND2xp33_ASAP7_75t_R n_7268 (.A(n_7266_o_0),
    .B(n_7267_o_0),
    .Y(n_7268_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7269 (.A1(n_7216_o_0),
    .A2(n_7196_o_0),
    .B(n_7232_o_0),
    .C(n_7219_o_0),
    .Y(n_7269_o_0));
 NAND4xp25_ASAP7_75t_R n_7270 (.A(n_7265_o_0),
    .B(n_7268_o_0),
    .C(n_7229_o_0),
    .D(n_7269_o_0),
    .Y(n_7270_o_0));
 OAI31xp33_ASAP7_75t_R n_7271 (.A1(n_7196_o_0),
    .A2(n_7202_o_0),
    .A3(n_7219_o_0),
    .B(n_7213_o_0),
    .Y(n_7271_o_0));
 INVx1_ASAP7_75t_R n_7272 (.A(n_7271_o_0),
    .Y(n_7272_o_0));
 OAI31xp33_ASAP7_75t_R n_7273 (.A1(n_7201_o_0),
    .A2(net46),
    .A3(n_7205_o_0),
    .B(n_7272_o_0),
    .Y(n_7273_o_0));
 OAI21xp33_ASAP7_75t_R n_7274 (.A1(n_7126_o_0),
    .A2(n_964_o_0),
    .B(n_7127_o_0),
    .Y(n_7274_o_0));
 INVx1_ASAP7_75t_R n_7275 (.A(n_7274_o_0),
    .Y(n_7275_o_0));
 AOI31xp33_ASAP7_75t_R n_7276 (.A1(n_7261_o_0),
    .A2(n_7270_o_0),
    .A3(n_7273_o_0),
    .B(n_7275_o_0),
    .Y(n_7276_o_0));
 OAI21xp33_ASAP7_75t_R n_7277 (.A1(n_7134_o_0),
    .A2(n_7258_o_0),
    .B(n_7276_o_0),
    .Y(n_7277_o_0));
 OAI21xp33_ASAP7_75t_R n_7278 (.A1(n_7127_o_1),
    .A2(n_7248_o_0),
    .B(n_7277_o_0),
    .Y(n_7278_o_0));
 INVx1_ASAP7_75t_R n_7279 (.A(n_7134_o_0),
    .Y(n_7279_o_0));
 AOI21xp33_ASAP7_75t_R n_7280 (.A1(n_7179_o_0),
    .A2(n_7199_o_0),
    .B(n_7200_o_0),
    .Y(n_7280_o_0));
 NOR2xp33_ASAP7_75t_R n_7281 (.A(n_7179_o_0),
    .B(n_7196_o_0),
    .Y(n_7281_o_0));
 OR4x1_ASAP7_75t_R n_7282 (.A(n_7280_o_0),
    .B(n_7281_o_0),
    .C(n_7205_o_0),
    .D(n_7224_o_0),
    .Y(n_7282_o_0));
 NOR2xp33_ASAP7_75t_R n_7283 (.A(n_7200_o_0),
    .B(n_7199_o_0),
    .Y(n_7283_o_0));
 INVx1_ASAP7_75t_R n_7284 (.A(n_7283_o_0),
    .Y(n_7284_o_0));
 NAND3xp33_ASAP7_75t_R n_7285 (.A(n_7199_o_0),
    .B(n_7182_o_0),
    .C(n_7200_o_0),
    .Y(n_7285_o_0));
 NAND3xp33_ASAP7_75t_R n_7286 (.A(n_7284_o_0),
    .B(n_7285_o_0),
    .C(n_7205_o_0),
    .Y(n_7286_o_0));
 AOI21xp33_ASAP7_75t_R n_7287 (.A1(n_7282_o_0),
    .A2(n_7286_o_0),
    .B(n_7240_o_0),
    .Y(n_7287_o_0));
 NOR3xp33_ASAP7_75t_R n_7288 (.A(n_7201_o_0),
    .B(n_7182_o_0),
    .C(n_7200_o_0),
    .Y(n_7288_o_0));
 AOI211xp5_ASAP7_75t_R n_7289 (.A1(n_7200_o_0),
    .A2(n_7182_o_0),
    .B(n_7288_o_0),
    .C(n_7205_o_0),
    .Y(n_7289_o_0));
 INVx1_ASAP7_75t_R n_7290 (.A(n_7289_o_0),
    .Y(n_7290_o_0));
 NOR2xp33_ASAP7_75t_R n_7291 (.A(n_7196_o_0),
    .B(n_7199_o_0),
    .Y(n_7291_o_0));
 NOR2xp33_ASAP7_75t_R n_7292 (.A(n_7200_o_0),
    .B(n_7216_o_0),
    .Y(n_7292_o_0));
 OAI21xp33_ASAP7_75t_R n_7293 (.A1(n_7291_o_0),
    .A2(n_7292_o_0),
    .B(n_7224_o_0),
    .Y(n_7293_o_0));
 AOI21xp33_ASAP7_75t_R n_7294 (.A1(n_7290_o_0),
    .A2(n_7293_o_0),
    .B(n_7241_o_0),
    .Y(n_7294_o_0));
 NAND2xp33_ASAP7_75t_R n_7295 (.A(n_7196_o_0),
    .B(n_7202_o_0),
    .Y(n_7295_o_0));
 AOI21xp33_ASAP7_75t_R n_7296 (.A1(n_7179_o_0),
    .A2(n_7199_o_0),
    .B(n_7196_o_0),
    .Y(n_7296_o_0));
 INVx1_ASAP7_75t_R n_7297 (.A(n_7296_o_0),
    .Y(n_7297_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7298 (.A1(n_7196_o_0),
    .A2(net79),
    .B(n_7182_o_0),
    .C(n_7219_o_0),
    .Y(n_7298_o_0));
 AOI31xp33_ASAP7_75t_R n_7299 (.A1(n_7151_o_0),
    .A2(n_7295_o_0),
    .A3(n_7297_o_0),
    .B(n_7298_o_0),
    .Y(n_7299_o_0));
 NOR2xp33_ASAP7_75t_R n_7300 (.A(n_7179_o_0),
    .B(n_7201_o_0),
    .Y(n_7300_o_0));
 OAI21xp33_ASAP7_75t_R n_7301 (.A1(n_7200_o_0),
    .A2(n_7262_o_0),
    .B(n_7219_o_0),
    .Y(n_7301_o_0));
 AOI211xp5_ASAP7_75t_R n_7302 (.A1(n_7300_o_0),
    .A2(n_7200_o_0),
    .B(n_7301_o_0),
    .C(n_7240_o_0),
    .Y(n_7302_o_0));
 NAND2xp33_ASAP7_75t_R n_7303 (.A(n_7182_o_0),
    .B(net79),
    .Y(n_7303_o_0));
 NAND2xp33_ASAP7_75t_R n_7304 (.A(n_7182_o_0),
    .B(n_7199_o_0),
    .Y(n_7304_o_0));
 AOI21xp33_ASAP7_75t_R n_7305 (.A1(n_7196_o_0),
    .A2(n_7304_o_0),
    .B(n_7205_o_0),
    .Y(n_7305_o_0));
 OAI21xp33_ASAP7_75t_R n_7306 (.A1(n_7179_o_0),
    .A2(n_7196_o_0),
    .B(n_7224_o_0),
    .Y(n_7306_o_0));
 NOR2xp33_ASAP7_75t_R n_7307 (.A(n_7306_o_0),
    .B(n_7241_o_0),
    .Y(n_7307_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7308 (.A1(n_7303_o_0),
    .A2(n_7196_o_0),
    .B(n_7305_o_0),
    .C(n_7307_o_0),
    .Y(n_7308_o_0));
 OAI221xp5_ASAP7_75t_R n_7309 (.A1(n_7240_o_0),
    .A2(n_7299_o_0),
    .B1(n_7302_o_0),
    .B2(n_7308_o_0),
    .C(n_7279_o_0),
    .Y(n_7309_o_0));
 OAI31xp33_ASAP7_75t_R n_7310 (.A1(n_7279_o_0),
    .A2(n_7287_o_0),
    .A3(n_7294_o_0),
    .B(n_7309_o_0),
    .Y(n_7310_o_0));
 NOR2xp33_ASAP7_75t_R n_7311 (.A(n_7196_o_0),
    .B(n_7220_o_0),
    .Y(n_7311_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7312 (.A1(n_7192_o_0),
    .A2(n_7191_o_0),
    .B(n_7195_o_0),
    .C(n_7199_o_0),
    .Y(n_7312_o_0));
 OAI311xp33_ASAP7_75t_R n_7313 (.A1(n_7196_o_0),
    .A2(n_7223_o_0),
    .A3(n_7222_o_0),
    .B1(n_7205_o_0),
    .C1(n_7312_o_0),
    .Y(n_7313_o_0));
 OAI31xp33_ASAP7_75t_R n_7314 (.A1(n_7224_o_0),
    .A2(n_7250_o_0),
    .A3(n_7311_o_0),
    .B(n_7313_o_0),
    .Y(n_7314_o_0));
 OAI21xp33_ASAP7_75t_R n_7315 (.A1(n_7241_o_0),
    .A2(n_7314_o_0),
    .B(n_7260_o_0),
    .Y(n_7315_o_0));
 OAI21xp33_ASAP7_75t_R n_7316 (.A1(n_7179_o_0),
    .A2(n_7199_o_0),
    .B(n_7200_o_0),
    .Y(n_7316_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7317 (.A1(net46),
    .A2(n_7216_o_0),
    .B(n_7316_o_0),
    .C(n_7151_o_0),
    .Y(n_7317_o_0));
 NOR3xp33_ASAP7_75t_R n_7318 (.A(n_7317_o_0),
    .B(n_7305_o_0),
    .C(n_7240_o_0),
    .Y(n_7318_o_0));
 NAND4xp25_ASAP7_75t_R n_7319 (.A(n_7196_o_0),
    .B(n_7224_o_0),
    .C(n_7201_o_0),
    .D(n_7179_o_0),
    .Y(n_7319_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7320 (.A1(n_7183_o_0),
    .A2(n_7180_o_0),
    .B(n_7200_o_0),
    .C(n_7219_o_0),
    .Y(n_7320_o_0));
 AOI21xp33_ASAP7_75t_R n_7321 (.A1(n_7319_o_0),
    .A2(n_7320_o_0),
    .B(n_7229_o_0),
    .Y(n_7321_o_0));
 NOR3xp33_ASAP7_75t_R n_7322 (.A(n_7304_o_0),
    .B(n_7151_o_0),
    .C(n_7196_o_0),
    .Y(n_7322_o_0));
 AOI211xp5_ASAP7_75t_R n_7323 (.A1(n_7289_o_0),
    .A2(n_7240_o_0),
    .B(n_7321_o_0),
    .C(n_7322_o_0),
    .Y(n_7323_o_0));
 OAI22xp33_ASAP7_75t_R n_7324 (.A1(n_7315_o_0),
    .A2(n_7318_o_0),
    .B1(n_7260_o_0),
    .B2(n_7323_o_0),
    .Y(n_7324_o_0));
 NAND2xp33_ASAP7_75t_R n_7325 (.A(n_923_o_0),
    .B(n_7119_o_0),
    .Y(n_7325_o_0));
 OAI21xp33_ASAP7_75t_R n_7326 (.A1(n_7119_o_0),
    .A2(n_923_o_0),
    .B(n_7325_o_0),
    .Y(n_7326_o_0));
 INVx1_ASAP7_75t_R n_7327 (.A(n_7326_o_0),
    .Y(n_7327_o_0));
 AOI21xp33_ASAP7_75t_R n_7328 (.A1(n_7127_o_1),
    .A2(n_7324_o_0),
    .B(n_7327_o_0),
    .Y(n_7328_o_0));
 OA21x2_ASAP7_75t_R n_7329 (.A1(n_7274_o_0),
    .A2(n_7310_o_0),
    .B(n_7328_o_0),
    .Y(n_7329_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7330 (.A1(_00978_),
    .A2(n_7119_o_0),
    .B(n_7120_o_0),
    .C(n_7278_o_0),
    .D(n_7329_o_0),
    .Y(n_7330_o_0));
 OAI31xp33_ASAP7_75t_R n_7331 (.A1(n_7182_o_0),
    .A2(n_7196_o_0),
    .A3(n_7219_o_0),
    .B(n_7213_o_0),
    .Y(n_7331_o_0));
 NOR3xp33_ASAP7_75t_R n_7332 (.A(n_7216_o_0),
    .B(net46),
    .C(n_7219_o_0),
    .Y(n_7332_o_0));
 NOR2xp33_ASAP7_75t_R n_7333 (.A(net46),
    .B(n_7224_o_0),
    .Y(n_7333_o_0));
 NOR3xp33_ASAP7_75t_R n_7334 (.A(n_7202_o_0),
    .B(n_7196_o_0),
    .C(n_7224_o_0),
    .Y(n_7334_o_0));
 AO21x1_ASAP7_75t_R n_7335 (.A1(n_7216_o_0),
    .A2(n_7333_o_0),
    .B(n_7334_o_0),
    .Y(n_7335_o_0));
 NOR2xp33_ASAP7_75t_R n_7336 (.A(n_7196_o_0),
    .B(n_7216_o_0),
    .Y(n_7336_o_0));
 NOR2xp33_ASAP7_75t_R n_7337 (.A(n_7182_o_0),
    .B(n_7200_o_0),
    .Y(n_7337_o_0));
 OAI21xp33_ASAP7_75t_R n_7338 (.A1(n_7196_o_0),
    .A2(n_7199_o_0),
    .B(n_7151_o_0),
    .Y(n_7338_o_0));
 INVx1_ASAP7_75t_R n_7339 (.A(n_7338_o_0),
    .Y(n_7339_o_0));
 NAND2xp33_ASAP7_75t_R n_7340 (.A(n_7196_o_0),
    .B(n_7304_o_0),
    .Y(n_7340_o_0));
 AOI21xp33_ASAP7_75t_R n_7341 (.A1(n_7339_o_0),
    .A2(n_7340_o_0),
    .B(n_7241_o_0),
    .Y(n_7341_o_0));
 OAI31xp33_ASAP7_75t_R n_7342 (.A1(n_7219_o_0),
    .A2(n_7336_o_0),
    .A3(n_7337_o_0),
    .B(n_7341_o_0),
    .Y(n_7342_o_0));
 OAI31xp33_ASAP7_75t_R n_7343 (.A1(n_7331_o_0),
    .A2(n_7332_o_0),
    .A3(n_7335_o_0),
    .B(n_7342_o_0),
    .Y(n_7343_o_0));
 NOR2xp33_ASAP7_75t_R n_7344 (.A(n_7182_o_0),
    .B(n_7201_o_0),
    .Y(n_7344_o_0));
 OAI21xp33_ASAP7_75t_R n_7345 (.A1(n_7200_o_0),
    .A2(n_7344_o_0),
    .B(n_7224_o_0),
    .Y(n_7345_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7346 (.A1(n_7216_o_0),
    .A2(net46),
    .B(n_7345_o_0),
    .C(n_7241_o_0),
    .Y(n_7346_o_0));
 INVx1_ASAP7_75t_R n_7347 (.A(n_7202_o_0),
    .Y(n_7347_o_0));
 AOI211xp5_ASAP7_75t_R n_7348 (.A1(n_7347_o_0),
    .A2(n_7196_o_0),
    .B(n_7205_o_0),
    .C(n_7243_o_0),
    .Y(n_7348_o_0));
 OAI211xp5_ASAP7_75t_R n_7349 (.A1(n_7306_o_0),
    .A2(n_7288_o_0),
    .B(n_7320_o_0),
    .C(n_7229_o_0),
    .Y(n_7349_o_0));
 OAI211xp5_ASAP7_75t_R n_7350 (.A1(n_7346_o_0),
    .A2(n_7348_o_0),
    .B(n_7261_o_0),
    .C(n_7349_o_0),
    .Y(n_7350_o_0));
 OAI21xp33_ASAP7_75t_R n_7351 (.A1(n_7261_o_0),
    .A2(n_7343_o_0),
    .B(n_7350_o_0),
    .Y(n_7351_o_0));
 OAI21xp33_ASAP7_75t_R n_7352 (.A1(n_7196_o_0),
    .A2(n_7216_o_0),
    .B(n_7205_o_0),
    .Y(n_7352_o_0));
 NAND2xp33_ASAP7_75t_R n_7353 (.A(n_7182_o_0),
    .B(n_7199_o_0),
    .Y(n_7353_o_0));
 NAND3xp33_ASAP7_75t_R n_7354 (.A(n_7353_o_0),
    .B(n_7151_o_0),
    .C(net46),
    .Y(n_7354_o_0));
 OAI211xp5_ASAP7_75t_R n_7355 (.A1(net23),
    .A2(n_7352_o_0),
    .B(n_7354_o_0),
    .C(n_7279_o_0),
    .Y(n_7355_o_0));
 AOI211xp5_ASAP7_75t_R n_7356 (.A1(n_7179_o_0),
    .A2(net79),
    .B(n_7205_o_0),
    .C(net46),
    .Y(n_7356_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7357 (.A1(n_7201_o_0),
    .A2(net46),
    .B(n_7301_o_0),
    .C(n_7134_o_0),
    .Y(n_7357_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7358 (.A1(n_7201_o_0),
    .A2(n_7200_o_0),
    .B(n_7250_o_0),
    .C(n_7224_o_0),
    .Y(n_7358_o_0));
 INVx1_ASAP7_75t_R n_7359 (.A(n_7358_o_0),
    .Y(n_7359_o_0));
 OAI22xp33_ASAP7_75t_R n_7360 (.A1(n_7355_o_0),
    .A2(n_7356_o_0),
    .B1(n_7357_o_0),
    .B2(n_7359_o_0),
    .Y(n_7360_o_0));
 NAND2xp33_ASAP7_75t_R n_7361 (.A(n_7200_o_0),
    .B(n_7201_o_0),
    .Y(n_7361_o_0));
 INVx1_ASAP7_75t_R n_7362 (.A(n_7361_o_0),
    .Y(n_7362_o_0));
 NOR3xp33_ASAP7_75t_R n_7363 (.A(n_7279_o_0),
    .B(n_7224_o_0),
    .C(n_7362_o_0),
    .Y(n_7363_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7364 (.A1(n_7201_o_0),
    .A2(n_7233_o_0),
    .B(n_7255_o_0),
    .C(n_7241_o_0),
    .Y(n_7364_o_0));
 INVx1_ASAP7_75t_R n_7365 (.A(n_7364_o_0),
    .Y(n_7365_o_0));
 AOI21xp33_ASAP7_75t_R n_7366 (.A1(_00978_),
    .A2(n_7119_o_0),
    .B(n_7120_o_0),
    .Y(n_7366_o_0));
 INVx1_ASAP7_75t_R n_7367 (.A(n_7366_o_0),
    .Y(n_7367_o_0));
 OAI21xp33_ASAP7_75t_R n_7368 (.A1(n_7363_o_0),
    .A2(n_7365_o_0),
    .B(n_7367_o_0),
    .Y(n_7368_o_0));
 AOI21xp33_ASAP7_75t_R n_7369 (.A1(n_7213_o_0),
    .A2(n_7360_o_0),
    .B(n_7368_o_0),
    .Y(n_7369_o_0));
 AOI21xp33_ASAP7_75t_R n_7370 (.A1(n_7326_o_0),
    .A2(n_7351_o_0),
    .B(n_7369_o_0),
    .Y(n_7370_o_0));
 NOR3xp33_ASAP7_75t_R n_7371 (.A(n_7304_o_0),
    .B(n_7151_o_0),
    .C(net46),
    .Y(n_7371_o_0));
 OAI21xp33_ASAP7_75t_R n_7372 (.A1(n_7196_o_0),
    .A2(n_7202_o_0),
    .B(n_7205_o_0),
    .Y(n_7372_o_0));
 NOR2xp33_ASAP7_75t_R n_7373 (.A(n_7182_o_0),
    .B(n_7201_o_0),
    .Y(n_7373_o_0));
 OAI21xp33_ASAP7_75t_R n_7374 (.A1(net23),
    .A2(n_7373_o_0),
    .B(n_7219_o_0),
    .Y(n_7374_o_0));
 OAI211xp5_ASAP7_75t_R n_7375 (.A1(n_7372_o_0),
    .A2(n_7250_o_0),
    .B(n_7374_o_0),
    .C(n_7261_o_0),
    .Y(n_7375_o_0));
 OAI31xp33_ASAP7_75t_R n_7376 (.A1(n_7261_o_0),
    .A2(n_7348_o_0),
    .A3(n_7371_o_0),
    .B(n_7375_o_0),
    .Y(n_7376_o_0));
 NAND2xp33_ASAP7_75t_R n_7377 (.A(n_7179_o_0),
    .B(n_7200_o_0),
    .Y(n_7377_o_0));
 NAND2xp33_ASAP7_75t_R n_7378 (.A(n_7196_o_0),
    .B(n_7216_o_0),
    .Y(n_7378_o_0));
 NOR3xp33_ASAP7_75t_R n_7379 (.A(n_7196_o_0),
    .B(n_7201_o_0),
    .C(n_7179_o_0),
    .Y(n_7379_o_0));
 AOI211xp5_ASAP7_75t_R n_7380 (.A1(n_7202_o_0),
    .A2(n_7196_o_0),
    .B(n_7379_o_0),
    .C(n_7224_o_0),
    .Y(n_7380_o_0));
 AOI31xp33_ASAP7_75t_R n_7381 (.A1(n_7205_o_0),
    .A2(n_7377_o_0),
    .A3(n_7378_o_0),
    .B(n_7380_o_0),
    .Y(n_7381_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7382 (.A1(n_7182_o_0),
    .A2(n_7201_o_0),
    .B(n_7200_o_0),
    .C(n_7205_o_0),
    .Y(n_7382_o_0));
 NAND2xp33_ASAP7_75t_R n_7383 (.A(net79),
    .B(n_7382_o_0),
    .Y(n_7383_o_0));
 AOI21xp33_ASAP7_75t_R n_7384 (.A1(n_7179_o_0),
    .A2(net79),
    .B(net46),
    .Y(n_7384_o_0));
 AOI21xp33_ASAP7_75t_R n_7385 (.A1(n_7224_o_0),
    .A2(n_7384_o_0),
    .B(n_7261_o_0),
    .Y(n_7385_o_0));
 AOI21xp33_ASAP7_75t_R n_7386 (.A1(n_7383_o_0),
    .A2(n_7385_o_0),
    .B(n_7229_o_0),
    .Y(n_7386_o_0));
 OAI21xp33_ASAP7_75t_R n_7387 (.A1(n_7279_o_0),
    .A2(n_7381_o_0),
    .B(n_7386_o_0),
    .Y(n_7387_o_0));
 OAI211xp5_ASAP7_75t_R n_7388 (.A1(n_7241_o_0),
    .A2(n_7376_o_0),
    .B(n_7387_o_0),
    .C(n_7326_o_0),
    .Y(n_7388_o_0));
 OAI21xp33_ASAP7_75t_R n_7389 (.A1(n_7201_o_0),
    .A2(n_7196_o_0),
    .B(n_7151_o_0),
    .Y(n_7389_o_0));
 NAND2xp33_ASAP7_75t_R n_7390 (.A(n_7389_o_0),
    .B(n_7213_o_0),
    .Y(n_7390_o_0));
 AOI21xp33_ASAP7_75t_R n_7391 (.A1(n_7200_o_0),
    .A2(n_7202_o_0),
    .B(n_7205_o_0),
    .Y(n_7391_o_0));
 OAI21xp33_ASAP7_75t_R n_7392 (.A1(n_7200_o_0),
    .A2(n_7344_o_0),
    .B(n_7391_o_0),
    .Y(n_7392_o_0));
 NAND3xp33_ASAP7_75t_R n_7393 (.A(n_7392_o_0),
    .B(n_7265_o_0),
    .C(n_7229_o_0),
    .Y(n_7393_o_0));
 OAI31xp33_ASAP7_75t_R n_7394 (.A1(n_7283_o_0),
    .A2(n_7322_o_0),
    .A3(n_7390_o_0),
    .B(n_7393_o_0),
    .Y(n_7394_o_0));
 INVx1_ASAP7_75t_R n_7395 (.A(n_7234_o_0),
    .Y(n_7395_o_0));
 NOR2xp33_ASAP7_75t_R n_7396 (.A(n_7200_o_0),
    .B(n_7201_o_0),
    .Y(n_7396_o_0));
 NAND3xp33_ASAP7_75t_R n_7397 (.A(n_7303_o_0),
    .B(net46),
    .C(n_7219_o_0),
    .Y(n_7397_o_0));
 OAI311xp33_ASAP7_75t_R n_7398 (.A1(n_7219_o_0),
    .A2(n_7395_o_0),
    .A3(n_7396_o_0),
    .B1(n_7229_o_0),
    .C1(n_7397_o_0),
    .Y(n_7398_o_0));
 NOR2xp33_ASAP7_75t_R n_7399 (.A(n_7182_o_0),
    .B(n_7196_o_0),
    .Y(n_7399_o_0));
 OAI21xp33_ASAP7_75t_R n_7400 (.A1(n_7200_o_0),
    .A2(n_7262_o_0),
    .B(n_7224_o_0),
    .Y(n_7400_o_0));
 NAND2xp33_ASAP7_75t_R n_7401 (.A(n_7182_o_0),
    .B(n_7200_o_0),
    .Y(n_7401_o_0));
 INVx1_ASAP7_75t_R n_7402 (.A(n_7401_o_0),
    .Y(n_7402_o_0));
 OA21x2_ASAP7_75t_R n_7403 (.A1(n_7320_o_0),
    .A2(n_7402_o_0),
    .B(n_7241_o_0),
    .Y(n_7403_o_0));
 OAI21xp33_ASAP7_75t_R n_7404 (.A1(n_7399_o_0),
    .A2(n_7400_o_0),
    .B(n_7403_o_0),
    .Y(n_7404_o_0));
 AOI31xp33_ASAP7_75t_R n_7405 (.A1(n_7398_o_0),
    .A2(n_7404_o_0),
    .A3(n_7279_o_0),
    .B(n_7366_o_0),
    .Y(n_7405_o_0));
 OAI21xp33_ASAP7_75t_R n_7406 (.A1(n_7260_o_0),
    .A2(n_7394_o_0),
    .B(n_7405_o_0),
    .Y(n_7406_o_0));
 AOI21xp33_ASAP7_75t_R n_7407 (.A1(n_7388_o_0),
    .A2(n_7406_o_0),
    .B(n_7275_o_0),
    .Y(n_7407_o_0));
 AOI21xp33_ASAP7_75t_R n_7408 (.A1(n_7275_o_0),
    .A2(n_7370_o_0),
    .B(n_7407_o_0),
    .Y(n_7408_o_0));
 NOR2xp33_ASAP7_75t_R n_7409 (.A(n_7200_o_0),
    .B(n_7220_o_0),
    .Y(n_7409_o_0));
 AOI21xp33_ASAP7_75t_R n_7410 (.A1(n_7200_o_0),
    .A2(n_7344_o_0),
    .B(n_7219_o_0),
    .Y(n_7410_o_0));
 AOI21xp33_ASAP7_75t_R n_7411 (.A1(n_7233_o_0),
    .A2(n_7410_o_0),
    .B(n_7229_o_0),
    .Y(n_7411_o_0));
 OAI21xp33_ASAP7_75t_R n_7412 (.A1(n_7338_o_0),
    .A2(n_7409_o_0),
    .B(n_7411_o_0),
    .Y(n_7412_o_0));
 AOI211xp5_ASAP7_75t_R n_7413 (.A1(n_7182_o_0),
    .A2(n_7201_o_0),
    .B(n_7223_o_0),
    .C(n_7200_o_0),
    .Y(n_7413_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7414 (.A1(net79),
    .A2(net46),
    .B(n_7182_o_0),
    .C(n_7205_o_0),
    .D(n_7241_o_0),
    .Y(n_7414_o_0));
 OAI31xp33_ASAP7_75t_R n_7415 (.A1(n_7224_o_0),
    .A2(n_7197_o_0),
    .A3(n_7413_o_0),
    .B(n_7414_o_0),
    .Y(n_7415_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7416 (.A1(n_7344_o_0),
    .A2(n_7200_o_0),
    .B(n_7219_o_0),
    .C(n_7213_o_0),
    .Y(n_7416_o_0));
 INVx1_ASAP7_75t_R n_7417 (.A(n_7379_o_0),
    .Y(n_7417_o_0));
 AOI22xp33_ASAP7_75t_R n_7418 (.A1(n_7416_o_0),
    .A2(n_7319_o_0),
    .B1(n_7233_o_0),
    .B2(n_7417_o_0),
    .Y(n_7418_o_0));
 NAND3xp33_ASAP7_75t_R n_7419 (.A(n_7416_o_0),
    .B(n_7319_o_0),
    .C(n_7224_o_0),
    .Y(n_7419_o_0));
 NOR2xp33_ASAP7_75t_R n_7420 (.A(n_7201_o_0),
    .B(n_7224_o_0),
    .Y(n_7420_o_0));
 NAND3xp33_ASAP7_75t_R n_7421 (.A(n_7229_o_0),
    .B(n_7196_o_0),
    .C(n_7420_o_0),
    .Y(n_7421_o_0));
 OAI311xp33_ASAP7_75t_R n_7422 (.A1(n_7196_o_0),
    .A2(n_7213_o_0),
    .A3(n_7304_o_0),
    .B1(n_7261_o_0),
    .C1(n_7421_o_0),
    .Y(n_7422_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7423 (.A1(n_7224_o_0),
    .A2(n_7418_o_0),
    .B(n_7419_o_0),
    .C(n_7422_o_0),
    .Y(n_7423_o_0));
 AOI31xp33_ASAP7_75t_R n_7424 (.A1(n_7260_o_0),
    .A2(n_7412_o_0),
    .A3(n_7415_o_0),
    .B(n_7423_o_0),
    .Y(n_7424_o_0));
 AOI21xp33_ASAP7_75t_R n_7425 (.A1(n_7182_o_0),
    .A2(net79),
    .B(n_7196_o_0),
    .Y(n_7425_o_0));
 INVx1_ASAP7_75t_R n_7426 (.A(n_7251_o_0),
    .Y(n_7426_o_0));
 OAI21xp33_ASAP7_75t_R n_7427 (.A1(n_7425_o_0),
    .A2(n_7426_o_0),
    .B(n_7219_o_0),
    .Y(n_7427_o_0));
 OAI211xp5_ASAP7_75t_R n_7428 (.A1(n_7396_o_0),
    .A2(n_7372_o_0),
    .B(n_7427_o_0),
    .C(n_7229_o_0),
    .Y(n_7428_o_0));
 NOR2xp33_ASAP7_75t_R n_7429 (.A(n_7196_o_0),
    .B(n_7344_o_0),
    .Y(n_7429_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7430 (.A1(n_7179_o_0),
    .A2(net46),
    .B(n_7201_o_0),
    .C(n_7219_o_0),
    .Y(n_7430_o_0));
 OAI21xp33_ASAP7_75t_R n_7431 (.A1(n_7400_o_0),
    .A2(n_7429_o_0),
    .B(n_7430_o_0),
    .Y(n_7431_o_0));
 AOI21xp33_ASAP7_75t_R n_7432 (.A1(n_7241_o_0),
    .A2(n_7431_o_0),
    .B(n_7260_o_0),
    .Y(n_7432_o_0));
 AOI311xp33_ASAP7_75t_R n_7433 (.A1(n_7196_o_0),
    .A2(n_7180_o_0),
    .A3(n_7183_o_0),
    .B(n_7219_o_0),
    .C(n_7291_o_0),
    .Y(n_7433_o_0));
 INVx1_ASAP7_75t_R n_7434 (.A(n_7336_o_0),
    .Y(n_7434_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7435 (.A1(n_7151_o_0),
    .A2(n_7233_o_0),
    .B(n_7433_o_0),
    .C(n_7434_o_0),
    .Y(n_7435_o_0));
 NAND2xp33_ASAP7_75t_R n_7436 (.A(n_7205_o_0),
    .B(n_7285_o_0),
    .Y(n_7436_o_0));
 OAI221xp5_ASAP7_75t_R n_7437 (.A1(n_7201_o_0),
    .A2(n_7377_o_0),
    .B1(net46),
    .B2(n_7344_o_0),
    .C(n_7151_o_0),
    .Y(n_7437_o_0));
 NAND3xp33_ASAP7_75t_R n_7438 (.A(n_7436_o_0),
    .B(n_7437_o_0),
    .C(n_7240_o_0),
    .Y(n_7438_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7439 (.A1(n_7240_o_0),
    .A2(n_7435_o_0),
    .B(n_7438_o_0),
    .C(n_7134_o_0),
    .Y(n_7439_o_0));
 AOI211xp5_ASAP7_75t_R n_7440 (.A1(n_7428_o_0),
    .A2(n_7432_o_0),
    .B(n_7439_o_0),
    .C(n_7366_o_0),
    .Y(n_7440_o_0));
 AOI21xp33_ASAP7_75t_R n_7441 (.A1(n_7424_o_0),
    .A2(n_7326_o_0),
    .B(n_7440_o_0),
    .Y(n_7441_o_0));
 OAI21xp33_ASAP7_75t_R n_7442 (.A1(n_7303_o_0),
    .A2(net46),
    .B(n_7391_o_0),
    .Y(n_7442_o_0));
 OAI311xp33_ASAP7_75t_R n_7443 (.A1(n_7201_o_0),
    .A2(n_7151_o_0),
    .A3(net46),
    .B1(n_7229_o_0),
    .C1(n_7442_o_0),
    .Y(n_7443_o_0));
 OAI221xp5_ASAP7_75t_R n_7444 (.A1(net23),
    .A2(n_7338_o_0),
    .B1(n_7396_o_0),
    .B2(n_7372_o_0),
    .C(n_7241_o_0),
    .Y(n_7444_o_0));
 AND3x1_ASAP7_75t_R n_7445 (.A(n_7443_o_0),
    .B(n_7444_o_0),
    .C(n_7279_o_0),
    .Y(n_7445_o_0));
 INVx1_ASAP7_75t_R n_7446 (.A(n_7316_o_0),
    .Y(n_7446_o_0));
 OAI21xp33_ASAP7_75t_R n_7447 (.A1(n_7196_o_0),
    .A2(n_7202_o_0),
    .B(n_7219_o_0),
    .Y(n_7447_o_0));
 AO21x1_ASAP7_75t_R n_7448 (.A1(n_7196_o_0),
    .A2(n_7220_o_0),
    .B(n_7447_o_0),
    .Y(n_7448_o_0));
 OAI31xp33_ASAP7_75t_R n_7449 (.A1(n_7219_o_0),
    .A2(n_7446_o_0),
    .A3(n_7396_o_0),
    .B(n_7448_o_0),
    .Y(n_7449_o_0));
 OAI21xp33_ASAP7_75t_R n_7450 (.A1(n_7179_o_0),
    .A2(n_7199_o_0),
    .B(n_7219_o_0),
    .Y(n_7450_o_0));
 OAI21xp33_ASAP7_75t_R n_7451 (.A1(n_7263_o_0),
    .A2(n_7450_o_0),
    .B(n_7229_o_0),
    .Y(n_7451_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7452 (.A1(n_7205_o_0),
    .A2(n_7361_o_0),
    .B(n_7451_o_0),
    .C(n_7261_o_0),
    .Y(n_7452_o_0));
 AOI21xp33_ASAP7_75t_R n_7453 (.A1(n_7241_o_0),
    .A2(n_7449_o_0),
    .B(n_7452_o_0),
    .Y(n_7453_o_0));
 INVx1_ASAP7_75t_R n_7454 (.A(n_7225_o_0),
    .Y(n_7454_o_0));
 OAI21xp33_ASAP7_75t_R n_7455 (.A1(n_7425_o_0),
    .A2(n_7454_o_0),
    .B(n_7240_o_0),
    .Y(n_7455_o_0));
 NOR2xp33_ASAP7_75t_R n_7456 (.A(n_7201_o_0),
    .B(n_7233_o_0),
    .Y(n_7456_o_0));
 AOI21xp33_ASAP7_75t_R n_7457 (.A1(n_7179_o_0),
    .A2(n_7196_o_0),
    .B(n_7224_o_0),
    .Y(n_7457_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7458 (.A1(n_7201_o_0),
    .A2(n_7377_o_0),
    .B(n_7457_o_0),
    .C(n_7229_o_0),
    .Y(n_7458_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7459 (.A1(n_7456_o_0),
    .A2(n_7254_o_0),
    .B(n_7458_o_0),
    .C(n_7261_o_0),
    .Y(n_7459_o_0));
 OAI21xp33_ASAP7_75t_R n_7460 (.A1(n_7455_o_0),
    .A2(n_7218_o_0),
    .B(n_7459_o_0),
    .Y(n_7460_o_0));
 OAI21xp33_ASAP7_75t_R n_7461 (.A1(n_7200_o_0),
    .A2(n_7201_o_0),
    .B(n_7151_o_0),
    .Y(n_7461_o_0));
 NAND2xp33_ASAP7_75t_R n_7462 (.A(n_7461_o_0),
    .B(n_7436_o_0),
    .Y(n_7462_o_0));
 AOI31xp33_ASAP7_75t_R n_7463 (.A1(net79),
    .A2(net46),
    .A3(n_7224_o_0),
    .B(n_7240_o_0),
    .Y(n_7463_o_0));
 AOI21xp33_ASAP7_75t_R n_7464 (.A1(n_7430_o_0),
    .A2(n_7463_o_0),
    .B(n_7260_o_0),
    .Y(n_7464_o_0));
 OAI21xp33_ASAP7_75t_R n_7465 (.A1(n_7213_o_0),
    .A2(n_7462_o_0),
    .B(n_7464_o_0),
    .Y(n_7465_o_0));
 NAND3xp33_ASAP7_75t_R n_7466 (.A(n_7460_o_0),
    .B(n_7465_o_0),
    .C(n_7327_o_0),
    .Y(n_7466_o_0));
 OAI311xp33_ASAP7_75t_R n_7467 (.A1(n_7327_o_0),
    .A2(n_7445_o_0),
    .A3(n_7453_o_0),
    .B1(n_7127_o_1),
    .C1(n_7466_o_0),
    .Y(n_7467_o_0));
 OAI21xp33_ASAP7_75t_R n_7468 (.A1(n_7127_o_1),
    .A2(n_7441_o_0),
    .B(n_7467_o_0),
    .Y(n_7468_o_0));
 NAND2xp33_ASAP7_75t_R n_7469 (.A(n_7312_o_0),
    .B(n_7255_o_0),
    .Y(n_7469_o_0));
 OAI21xp33_ASAP7_75t_R n_7470 (.A1(n_7197_o_0),
    .A2(n_7292_o_0),
    .B(n_7219_o_0),
    .Y(n_7470_o_0));
 INVx1_ASAP7_75t_R n_7471 (.A(n_7242_o_0),
    .Y(n_7471_o_0));
 OAI21xp33_ASAP7_75t_R n_7472 (.A1(n_7200_o_0),
    .A2(n_7182_o_0),
    .B(n_7151_o_0),
    .Y(n_7472_o_0));
 OAI21xp33_ASAP7_75t_R n_7473 (.A1(n_7472_o_0),
    .A2(n_7296_o_0),
    .B(n_7240_o_0),
    .Y(n_7473_o_0));
 AOI21xp33_ASAP7_75t_R n_7474 (.A1(n_7401_o_0),
    .A2(n_7471_o_0),
    .B(n_7473_o_0),
    .Y(n_7474_o_0));
 AOI31xp33_ASAP7_75t_R n_7475 (.A1(n_7241_o_0),
    .A2(n_7469_o_0),
    .A3(n_7470_o_0),
    .B(n_7474_o_0),
    .Y(n_7475_o_0));
 AOI211xp5_ASAP7_75t_R n_7476 (.A1(n_7183_o_0),
    .A2(n_7180_o_0),
    .B(n_7151_o_0),
    .C(n_7200_o_0),
    .Y(n_7476_o_0));
 AOI21xp33_ASAP7_75t_R n_7477 (.A1(n_7219_o_0),
    .A2(n_7292_o_0),
    .B(n_7476_o_0),
    .Y(n_7477_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7478 (.A1(n_7224_o_0),
    .A2(n_7409_o_0),
    .B(n_7414_o_0),
    .C(n_7261_o_0),
    .Y(n_7478_o_0));
 OAI21xp33_ASAP7_75t_R n_7479 (.A1(n_7229_o_0),
    .A2(n_7477_o_0),
    .B(n_7478_o_0),
    .Y(n_7479_o_0));
 OAI21xp33_ASAP7_75t_R n_7480 (.A1(n_7279_o_0),
    .A2(n_7475_o_0),
    .B(n_7479_o_0),
    .Y(n_7480_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7481 (.A1(n_7196_o_0),
    .A2(net79),
    .B(n_7179_o_0),
    .C(n_7219_o_0),
    .Y(n_7481_o_0));
 AOI21xp33_ASAP7_75t_R n_7482 (.A1(n_7179_o_0),
    .A2(n_7201_o_0),
    .B(n_7196_o_0),
    .Y(n_7482_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7483 (.A1(n_7472_o_0),
    .A2(n_7482_o_0),
    .B(n_7364_o_0),
    .C(n_7279_o_0),
    .Y(n_7483_o_0));
 NAND2xp33_ASAP7_75t_R n_7484 (.A(n_7241_o_0),
    .B(n_7481_o_0),
    .Y(n_7484_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7485 (.A1(n_7196_o_0),
    .A2(n_7221_o_0),
    .B(n_7281_o_0),
    .C(n_7219_o_0),
    .D(n_7240_o_0),
    .Y(n_7485_o_0));
 OAI21xp33_ASAP7_75t_R n_7486 (.A1(n_7242_o_0),
    .A2(n_7429_o_0),
    .B(n_7485_o_0),
    .Y(n_7486_o_0));
 OAI311xp33_ASAP7_75t_R n_7487 (.A1(n_7219_o_0),
    .A2(n_7395_o_0),
    .A3(n_7396_o_0),
    .B1(n_7229_o_0),
    .C1(n_7269_o_0),
    .Y(n_7487_o_0));
 AO31x2_ASAP7_75t_R n_7488 (.A1(n_7486_o_0),
    .A2(n_7487_o_0),
    .A3(n_7279_o_0),
    .B(n_7327_o_0),
    .Y(n_7488_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7489 (.A1(n_7241_o_0),
    .A2(n_7481_o_0),
    .B(n_7483_o_0),
    .C(n_7484_o_0),
    .D(n_7488_o_0),
    .Y(n_7489_o_0));
 AOI21xp33_ASAP7_75t_R n_7490 (.A1(n_7367_o_0),
    .A2(n_7480_o_0),
    .B(n_7489_o_0),
    .Y(n_7490_o_0));
 NOR2xp33_ASAP7_75t_R n_7491 (.A(n_7244_o_0),
    .B(n_7338_o_0),
    .Y(n_7491_o_0));
 NOR2xp33_ASAP7_75t_R n_7492 (.A(n_7384_o_0),
    .B(n_7372_o_0),
    .Y(n_7492_o_0));
 AOI211xp5_ASAP7_75t_R n_7493 (.A1(n_7491_o_0),
    .A2(n_7377_o_0),
    .B(n_7492_o_0),
    .C(n_7241_o_0),
    .Y(n_7493_o_0));
 AOI21xp33_ASAP7_75t_R n_7494 (.A1(net46),
    .A2(n_7220_o_0),
    .B(n_7242_o_0),
    .Y(n_7494_o_0));
 NOR3xp33_ASAP7_75t_R n_7495 (.A(n_7399_o_0),
    .B(n_7300_o_0),
    .C(n_7205_o_0),
    .Y(n_7495_o_0));
 NOR3xp33_ASAP7_75t_R n_7496 (.A(n_7494_o_0),
    .B(n_7495_o_0),
    .C(n_7240_o_0),
    .Y(n_7496_o_0));
 INVx1_ASAP7_75t_R n_7497 (.A(n_7482_o_0),
    .Y(n_7497_o_0));
 OAI211xp5_ASAP7_75t_R n_7498 (.A1(n_7202_o_0),
    .A2(net46),
    .B(n_7497_o_0),
    .C(n_7205_o_0),
    .Y(n_7498_o_0));
 OAI21xp33_ASAP7_75t_R n_7499 (.A1(n_7337_o_0),
    .A2(n_7231_o_0),
    .B(n_7224_o_0),
    .Y(n_7499_o_0));
 AOI31xp33_ASAP7_75t_R n_7500 (.A1(n_7229_o_0),
    .A2(n_7499_o_0),
    .A3(n_7285_o_0),
    .B(n_7260_o_0),
    .Y(n_7500_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7501 (.A1(n_7498_o_0),
    .A2(n_7383_o_0),
    .B(n_7229_o_0),
    .C(n_7500_o_0),
    .Y(n_7501_o_0));
 OAI31xp33_ASAP7_75t_R n_7502 (.A1(n_7261_o_0),
    .A2(n_7493_o_0),
    .A3(n_7496_o_0),
    .B(n_7501_o_0),
    .Y(n_7502_o_0));
 NOR3xp33_ASAP7_75t_R n_7503 (.A(n_7232_o_0),
    .B(n_7244_o_0),
    .C(n_7219_o_0),
    .Y(n_7503_o_0));
 NOR2xp33_ASAP7_75t_R n_7504 (.A(n_7200_o_0),
    .B(n_7266_o_0),
    .Y(n_7504_o_0));
 OAI31xp33_ASAP7_75t_R n_7505 (.A1(n_7224_o_0),
    .A2(n_7504_o_0),
    .A3(n_7197_o_0),
    .B(n_7213_o_0),
    .Y(n_7505_o_0));
 NAND2xp33_ASAP7_75t_R n_7506 (.A(n_7200_o_0),
    .B(n_7201_o_0),
    .Y(n_7506_o_0));
 OAI311xp33_ASAP7_75t_R n_7507 (.A1(net46),
    .A2(n_7223_o_0),
    .A3(n_7222_o_0),
    .B1(n_7205_o_0),
    .C1(n_7506_o_0),
    .Y(n_7507_o_0));
 OAI31xp33_ASAP7_75t_R n_7508 (.A1(n_7224_o_0),
    .A2(n_7280_o_0),
    .A3(n_7425_o_0),
    .B(n_7507_o_0),
    .Y(n_7508_o_0));
 AOI21xp33_ASAP7_75t_R n_7509 (.A1(n_7229_o_0),
    .A2(n_7508_o_0),
    .B(n_7261_o_0),
    .Y(n_7509_o_0));
 OAI21xp33_ASAP7_75t_R n_7510 (.A1(n_7503_o_0),
    .A2(n_7505_o_0),
    .B(n_7509_o_0),
    .Y(n_7510_o_0));
 OAI32xp33_ASAP7_75t_R n_7511 (.A1(n_7219_o_0),
    .A2(n_7291_o_0),
    .A3(n_7250_o_0),
    .B1(n_7197_o_0),
    .B2(n_7224_o_0),
    .Y(n_7511_o_0));
 INVx1_ASAP7_75t_R n_7512 (.A(n_7511_o_0),
    .Y(n_7512_o_0));
 OAI31xp33_ASAP7_75t_R n_7513 (.A1(n_7219_o_0),
    .A2(n_7231_o_0),
    .A3(n_7337_o_0),
    .B(n_7240_o_0),
    .Y(n_7513_o_0));
 AOI21xp33_ASAP7_75t_R n_7514 (.A1(n_7225_o_0),
    .A2(n_7506_o_0),
    .B(n_7513_o_0),
    .Y(n_7514_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7515 (.A1(n_7512_o_0),
    .A2(n_7213_o_0),
    .B(n_7514_o_0),
    .C(n_7261_o_0),
    .Y(n_7515_o_0));
 AOI31xp33_ASAP7_75t_R n_7516 (.A1(n_7327_o_0),
    .A2(n_7510_o_0),
    .A3(n_7515_o_0),
    .B(n_7275_o_0),
    .Y(n_7516_o_0));
 OAI21xp33_ASAP7_75t_R n_7517 (.A1(n_7367_o_0),
    .A2(n_7502_o_0),
    .B(n_7516_o_0),
    .Y(n_7517_o_0));
 OA21x2_ASAP7_75t_R n_7518 (.A1(n_7490_o_0),
    .A2(n_7127_o_1),
    .B(n_7517_o_0),
    .Y(n_7518_o_0));
 INVx1_ASAP7_75t_R n_7519 (.A(n_7127_o_1),
    .Y(n_7519_o_0));
 INVx1_ASAP7_75t_R n_7520 (.A(n_7400_o_0),
    .Y(n_7520_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7521 (.A1(n_7196_o_0),
    .A2(n_7202_o_0),
    .B(n_7520_o_0),
    .C(n_7261_o_0),
    .Y(n_7521_o_0));
 AOI21xp33_ASAP7_75t_R n_7522 (.A1(n_7182_o_0),
    .A2(n_7224_o_0),
    .B(net46),
    .Y(n_7522_o_0));
 AOI21xp33_ASAP7_75t_R n_7523 (.A1(n_7205_o_0),
    .A2(n_7429_o_0),
    .B(n_7522_o_0),
    .Y(n_7523_o_0));
 OAI21xp33_ASAP7_75t_R n_7524 (.A1(n_7279_o_0),
    .A2(n_7523_o_0),
    .B(n_7240_o_0),
    .Y(n_7524_o_0));
 AOI21xp33_ASAP7_75t_R n_7525 (.A1(n_7290_o_0),
    .A2(n_7521_o_0),
    .B(n_7524_o_0),
    .Y(n_7525_o_0));
 AOI21xp33_ASAP7_75t_R n_7526 (.A1(n_7506_o_0),
    .A2(n_7378_o_0),
    .B(n_7151_o_0),
    .Y(n_7526_o_0));
 AOI21xp33_ASAP7_75t_R n_7527 (.A1(n_7200_o_0),
    .A2(n_7216_o_0),
    .B(n_7151_o_0),
    .Y(n_7527_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7528 (.A1(n_7201_o_0),
    .A2(n_7377_o_0),
    .B(n_7151_o_0),
    .C(n_7527_o_0),
    .Y(n_7528_o_0));
 AOI21xp33_ASAP7_75t_R n_7529 (.A1(n_7260_o_0),
    .A2(n_7528_o_0),
    .B(n_7229_o_0),
    .Y(n_7529_o_0));
 OA21x2_ASAP7_75t_R n_7530 (.A1(n_7357_o_0),
    .A2(n_7526_o_0),
    .B(n_7529_o_0),
    .Y(n_7530_o_0));
 OAI211xp5_ASAP7_75t_R n_7531 (.A1(n_7219_o_0),
    .A2(n_7344_o_0),
    .B(n_7447_o_0),
    .C(n_7279_o_0),
    .Y(n_7531_o_0));
 OAI31xp33_ASAP7_75t_R n_7532 (.A1(n_7279_o_0),
    .A2(n_7317_o_0),
    .A3(n_7495_o_0),
    .B(n_7531_o_0),
    .Y(n_7532_o_0));
 NOR3xp33_ASAP7_75t_R n_7533 (.A(n_7311_o_0),
    .B(net23),
    .C(n_7224_o_0),
    .Y(n_7533_o_0));
 NOR3xp33_ASAP7_75t_R n_7534 (.A(n_7283_o_0),
    .B(n_7373_o_0),
    .C(n_7219_o_0),
    .Y(n_7534_o_0));
 OA21x2_ASAP7_75t_R n_7535 (.A1(n_7533_o_0),
    .A2(n_7534_o_0),
    .B(n_7134_o_0),
    .Y(n_7535_o_0));
 NAND2xp33_ASAP7_75t_R n_7536 (.A(n_7249_o_0),
    .B(n_7284_o_0),
    .Y(n_7536_o_0));
 OAI31xp33_ASAP7_75t_R n_7537 (.A1(net46),
    .A2(n_7219_o_0),
    .A3(n_7231_o_0),
    .B(n_7536_o_0),
    .Y(n_7537_o_0));
 OAI21xp33_ASAP7_75t_R n_7538 (.A1(n_7134_o_0),
    .A2(n_7537_o_0),
    .B(n_7241_o_0),
    .Y(n_7538_o_0));
 OAI221xp5_ASAP7_75t_R n_7539 (.A1(n_7241_o_0),
    .A2(n_7532_o_0),
    .B1(n_7535_o_0),
    .B2(n_7538_o_0),
    .C(n_7367_o_0),
    .Y(n_7539_o_0));
 OAI31xp33_ASAP7_75t_R n_7540 (.A1(n_7327_o_0),
    .A2(n_7525_o_0),
    .A3(n_7530_o_0),
    .B(n_7539_o_0),
    .Y(n_7540_o_0));
 INVx1_ASAP7_75t_R n_7541 (.A(n_7334_o_0),
    .Y(n_7541_o_0));
 AOI211xp5_ASAP7_75t_R n_7542 (.A1(n_7267_o_0),
    .A2(n_7262_o_0),
    .B(n_7409_o_0),
    .C(n_7240_o_0),
    .Y(n_7542_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7543 (.A1(n_7199_o_0),
    .A2(n_7179_o_0),
    .B(n_7200_o_0),
    .C(n_7205_o_0),
    .Y(n_7543_o_0));
 OAI21xp33_ASAP7_75t_R n_7544 (.A1(n_7197_o_0),
    .A2(n_7543_o_0),
    .B(n_7240_o_0),
    .Y(n_7544_o_0));
 AOI21xp33_ASAP7_75t_R n_7545 (.A1(n_7251_o_0),
    .A2(n_7249_o_0),
    .B(n_7544_o_0),
    .Y(n_7545_o_0));
 AOI21xp33_ASAP7_75t_R n_7546 (.A1(n_7541_o_0),
    .A2(n_7542_o_0),
    .B(n_7545_o_0),
    .Y(n_7546_o_0));
 OAI21xp33_ASAP7_75t_R n_7547 (.A1(n_7179_o_0),
    .A2(net46),
    .B(n_7229_o_0),
    .Y(n_7547_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7548 (.A1(n_7266_o_0),
    .A2(n_7196_o_0),
    .B(n_7249_o_0),
    .C(n_7241_o_0),
    .Y(n_7548_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7549 (.A1(n_7389_o_0),
    .A2(n_7352_o_0),
    .B(n_7547_o_0),
    .C(n_7548_o_0),
    .Y(n_7549_o_0));
 OAI22xp33_ASAP7_75t_R n_7550 (.A1(n_7546_o_0),
    .A2(n_7326_o_0),
    .B1(n_7367_o_0),
    .B2(n_7549_o_0),
    .Y(n_7550_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7551 (.A1(net79),
    .A2(net46),
    .B(n_7504_o_0),
    .C(n_7219_o_0),
    .Y(n_7551_o_0));
 AOI21xp33_ASAP7_75t_R n_7552 (.A1(n_7265_o_0),
    .A2(n_7551_o_0),
    .B(n_7241_o_0),
    .Y(n_7552_o_0));
 AOI21xp33_ASAP7_75t_R n_7553 (.A1(net79),
    .A2(n_7250_o_0),
    .B(n_7338_o_0),
    .Y(n_7553_o_0));
 AOI31xp33_ASAP7_75t_R n_7554 (.A1(n_7205_o_0),
    .A2(n_7340_o_0),
    .A3(n_7297_o_0),
    .B(n_7553_o_0),
    .Y(n_7554_o_0));
 OAI21xp33_ASAP7_75t_R n_7555 (.A1(n_7240_o_0),
    .A2(n_7554_o_0),
    .B(n_7327_o_0),
    .Y(n_7555_o_0));
 AOI21xp33_ASAP7_75t_R n_7556 (.A1(n_7506_o_0),
    .A2(n_7353_o_0),
    .B(n_7151_o_0),
    .Y(n_7556_o_0));
 AOI21xp33_ASAP7_75t_R n_7557 (.A1(n_7312_o_0),
    .A2(n_7316_o_0),
    .B(n_7205_o_0),
    .Y(n_7557_o_0));
 OAI211xp5_ASAP7_75t_R n_7558 (.A1(n_7450_o_0),
    .A2(n_7263_o_0),
    .B(n_7358_o_0),
    .C(n_7229_o_0),
    .Y(n_7558_o_0));
 OAI31xp33_ASAP7_75t_R n_7559 (.A1(n_7240_o_0),
    .A2(n_7556_o_0),
    .A3(n_7557_o_0),
    .B(n_7558_o_0),
    .Y(n_7559_o_0));
 AOI21xp33_ASAP7_75t_R n_7560 (.A1(n_7326_o_0),
    .A2(n_7559_o_0),
    .B(n_7260_o_0),
    .Y(n_7560_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7561 (.A1(n_7552_o_0),
    .A2(n_7555_o_0),
    .B(n_7560_o_0),
    .C(n_7275_o_0),
    .Y(n_7561_o_0));
 OA21x2_ASAP7_75t_R n_7562 (.A1(n_7134_o_0),
    .A2(n_7550_o_0),
    .B(n_7561_o_0),
    .Y(n_7562_o_0));
 AOI21xp33_ASAP7_75t_R n_7563 (.A1(n_7519_o_0),
    .A2(n_7540_o_0),
    .B(n_7562_o_0),
    .Y(n_7563_o_0));
 AOI211xp5_ASAP7_75t_R n_7564 (.A1(n_7210_o_0),
    .A2(net),
    .B(_00976_),
    .C(n_7211_o_0),
    .Y(n_7564_o_0));
 NAND3xp33_ASAP7_75t_R n_7565 (.A(n_7497_o_0),
    .B(n_7251_o_0),
    .C(n_7205_o_0),
    .Y(n_7565_o_0));
 OAI31xp33_ASAP7_75t_R n_7566 (.A1(n_7179_o_0),
    .A2(n_7224_o_0),
    .A3(n_7425_o_0),
    .B(n_7565_o_0),
    .Y(n_7566_o_0));
 OAI21xp33_ASAP7_75t_R n_7567 (.A1(n_7564_o_0),
    .A2(n_7239_o_0),
    .B(n_7566_o_0),
    .Y(n_7567_o_0));
 OAI211xp5_ASAP7_75t_R n_7568 (.A1(n_7196_o_0),
    .A2(n_7344_o_0),
    .B(n_7305_o_0),
    .C(n_7240_o_0),
    .Y(n_7568_o_0));
 OA21x2_ASAP7_75t_R n_7569 (.A1(n_7293_o_0),
    .A2(n_7241_o_0),
    .B(n_7260_o_0),
    .Y(n_7569_o_0));
 OAI21xp33_ASAP7_75t_R n_7570 (.A1(n_7281_o_0),
    .A2(n_7409_o_0),
    .B(n_7219_o_0),
    .Y(n_7570_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7571 (.A1(n_7180_o_0),
    .A2(n_7183_o_0),
    .B(net46),
    .C(n_7224_o_0),
    .D(n_7213_o_0),
    .Y(n_7571_o_0));
 AOI22xp33_ASAP7_75t_R n_7572 (.A1(n_7397_o_0),
    .A2(n_7400_o_0),
    .B1(n_7570_o_0),
    .B2(n_7571_o_0),
    .Y(n_7572_o_0));
 NAND3xp33_ASAP7_75t_R n_7573 (.A(n_7570_o_0),
    .B(n_7571_o_0),
    .C(n_7240_o_0),
    .Y(n_7573_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7574 (.A1(n_7240_o_0),
    .A2(n_7572_o_0),
    .B(n_7573_o_0),
    .C(n_7279_o_0),
    .Y(n_7574_o_0));
 AOI31xp33_ASAP7_75t_R n_7575 (.A1(n_7567_o_0),
    .A2(n_7568_o_0),
    .A3(n_7569_o_0),
    .B(n_7574_o_0),
    .Y(n_7575_o_0));
 OAI21xp33_ASAP7_75t_R n_7576 (.A1(n_7527_o_0),
    .A2(n_7334_o_0),
    .B(n_7312_o_0),
    .Y(n_7576_o_0));
 AOI21xp33_ASAP7_75t_R n_7577 (.A1(n_7225_o_0),
    .A2(n_7316_o_0),
    .B(n_7410_o_0),
    .Y(n_7577_o_0));
 AOI21xp33_ASAP7_75t_R n_7578 (.A1(n_7229_o_0),
    .A2(n_7577_o_0),
    .B(n_7260_o_0),
    .Y(n_7578_o_0));
 OAI21xp33_ASAP7_75t_R n_7579 (.A1(n_7240_o_0),
    .A2(n_7576_o_0),
    .B(n_7578_o_0),
    .Y(n_7579_o_0));
 OAI21xp33_ASAP7_75t_R n_7580 (.A1(n_7179_o_0),
    .A2(n_7196_o_0),
    .B(n_7205_o_0),
    .Y(n_7580_o_0));
 OAI21xp33_ASAP7_75t_R n_7581 (.A1(n_7373_o_0),
    .A2(n_7580_o_0),
    .B(n_7213_o_0),
    .Y(n_7581_o_0));
 NOR3xp33_ASAP7_75t_R n_7582 (.A(n_7384_o_0),
    .B(n_7482_o_0),
    .C(n_7224_o_0),
    .Y(n_7582_o_0));
 OAI21xp33_ASAP7_75t_R n_7583 (.A1(n_7420_o_0),
    .A2(n_7534_o_0),
    .B(n_7229_o_0),
    .Y(n_7583_o_0));
 OAI211xp5_ASAP7_75t_R n_7584 (.A1(n_7581_o_0),
    .A2(n_7582_o_0),
    .B(n_7583_o_0),
    .C(n_7260_o_0),
    .Y(n_7584_o_0));
 AO21x1_ASAP7_75t_R n_7585 (.A1(n_7579_o_0),
    .A2(n_7584_o_0),
    .B(n_7366_o_0),
    .Y(n_7585_o_0));
 OAI21xp33_ASAP7_75t_R n_7586 (.A1(n_7327_o_0),
    .A2(n_7575_o_0),
    .B(n_7585_o_0),
    .Y(n_7586_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7587 (.A1(n_7337_o_0),
    .A2(n_7322_o_0),
    .B(n_7224_o_0),
    .C(n_7289_o_0),
    .Y(n_7587_o_0));
 AOI31xp33_ASAP7_75t_R n_7588 (.A1(n_7205_o_0),
    .A2(n_7234_o_0),
    .A3(n_7233_o_0),
    .B(n_7134_o_0),
    .Y(n_7588_o_0));
 OA21x2_ASAP7_75t_R n_7589 (.A1(n_7182_o_0),
    .A2(n_7224_o_0),
    .B(n_7588_o_0),
    .Y(n_7589_o_0));
 AOI211xp5_ASAP7_75t_R n_7590 (.A1(n_7134_o_0),
    .A2(n_7587_o_0),
    .B(n_7589_o_0),
    .C(n_7213_o_0),
    .Y(n_7590_o_0));
 NOR2xp33_ASAP7_75t_R n_7591 (.A(n_7482_o_0),
    .B(n_7283_o_0),
    .Y(n_7591_o_0));
 AO22x1_ASAP7_75t_R n_7592 (.A1(n_7225_o_0),
    .A2(n_7285_o_0),
    .B1(n_7591_o_0),
    .B2(n_7205_o_0),
    .Y(n_7592_o_0));
 AOI21xp33_ASAP7_75t_R n_7593 (.A1(n_7219_o_0),
    .A2(n_7482_o_0),
    .B(n_7279_o_0),
    .Y(n_7593_o_0));
 OAI31xp33_ASAP7_75t_R n_7594 (.A1(n_7219_o_0),
    .A2(n_7296_o_0),
    .A3(n_7456_o_0),
    .B(n_7593_o_0),
    .Y(n_7594_o_0));
 OAI21xp33_ASAP7_75t_R n_7595 (.A1(n_7134_o_0),
    .A2(n_7592_o_0),
    .B(n_7594_o_0),
    .Y(n_7595_o_0));
 OAI21xp33_ASAP7_75t_R n_7596 (.A1(n_7229_o_0),
    .A2(n_7595_o_0),
    .B(n_7326_o_0),
    .Y(n_7596_o_0));
 OAI21xp33_ASAP7_75t_R n_7597 (.A1(n_7382_o_0),
    .A2(n_7322_o_0),
    .B(n_7279_o_0),
    .Y(n_7597_o_0));
 OAI21xp33_ASAP7_75t_R n_7598 (.A1(n_7196_o_0),
    .A2(n_7220_o_0),
    .B(n_7225_o_0),
    .Y(n_7598_o_0));
 OAI31xp33_ASAP7_75t_R n_7599 (.A1(n_7219_o_0),
    .A2(n_7296_o_0),
    .A3(n_7413_o_0),
    .B(n_7598_o_0),
    .Y(n_7599_o_0));
 AOI21xp33_ASAP7_75t_R n_7600 (.A1(n_7134_o_0),
    .A2(n_7599_o_0),
    .B(n_7229_o_0),
    .Y(n_7600_o_0));
 OAI22xp33_ASAP7_75t_R n_7601 (.A1(n_7456_o_0),
    .A2(n_7219_o_0),
    .B1(n_7221_o_0),
    .B2(n_7224_o_0),
    .Y(n_7601_o_0));
 AOI21xp33_ASAP7_75t_R n_7602 (.A1(n_7260_o_0),
    .A2(n_7457_o_0),
    .B(n_7241_o_0),
    .Y(n_7602_o_0));
 OAI21xp33_ASAP7_75t_R n_7603 (.A1(n_7456_o_0),
    .A2(n_7436_o_0),
    .B(n_7602_o_0),
    .Y(n_7603_o_0));
 AOI21xp33_ASAP7_75t_R n_7604 (.A1(n_7134_o_0),
    .A2(n_7601_o_0),
    .B(n_7603_o_0),
    .Y(n_7604_o_0));
 NAND2xp33_ASAP7_75t_R n_7605 (.A(n_7366_o_0),
    .B(n_7275_o_0),
    .Y(n_7605_o_0));
 AOI211xp5_ASAP7_75t_R n_7606 (.A1(n_7600_o_0),
    .A2(n_7597_o_0),
    .B(n_7604_o_0),
    .C(n_7275_o_0),
    .Y(n_7606_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7607 (.A1(n_7597_o_0),
    .A2(n_7600_o_0),
    .B(n_7604_o_0),
    .C(n_7605_o_0),
    .D(n_7606_o_0),
    .Y(n_7607_o_0));
 OAI21xp33_ASAP7_75t_R n_7608 (.A1(n_7590_o_0),
    .A2(n_7596_o_0),
    .B(n_7607_o_0),
    .Y(n_7608_o_0));
 OAI21xp33_ASAP7_75t_R n_7609 (.A1(n_7519_o_0),
    .A2(n_7586_o_0),
    .B(n_7608_o_0),
    .Y(n_7609_o_0));
 AOI211xp5_ASAP7_75t_R n_7610 (.A1(n_7436_o_0),
    .A2(n_7461_o_0),
    .B(n_7476_o_0),
    .C(n_7240_o_0),
    .Y(n_7610_o_0));
 INVx1_ASAP7_75t_R n_7611 (.A(n_7610_o_0),
    .Y(n_7611_o_0));
 INVx1_ASAP7_75t_R n_7612 (.A(n_7285_o_0),
    .Y(n_7612_o_0));
 INVx1_ASAP7_75t_R n_7613 (.A(n_7413_o_0),
    .Y(n_7613_o_0));
 NAND2xp33_ASAP7_75t_R n_7614 (.A(n_7527_o_0),
    .B(n_7613_o_0),
    .Y(n_7614_o_0));
 OAI31xp33_ASAP7_75t_R n_7615 (.A1(n_7224_o_0),
    .A2(n_7612_o_0),
    .A3(n_7283_o_0),
    .B(n_7614_o_0),
    .Y(n_7615_o_0));
 AOI21xp33_ASAP7_75t_R n_7616 (.A1(n_7229_o_0),
    .A2(n_7615_o_0),
    .B(n_7134_o_0),
    .Y(n_7616_o_0));
 NAND2xp33_ASAP7_75t_R n_7617 (.A(n_7179_o_0),
    .B(n_7196_o_0),
    .Y(n_7617_o_0));
 OAI211xp5_ASAP7_75t_R n_7618 (.A1(n_7202_o_0),
    .A2(n_7196_o_0),
    .B(n_7205_o_0),
    .C(n_7617_o_0),
    .Y(n_7618_o_0));
 OAI31xp33_ASAP7_75t_R n_7619 (.A1(n_7224_o_0),
    .A2(n_7426_o_0),
    .A3(n_7232_o_0),
    .B(n_7618_o_0),
    .Y(n_7619_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7620 (.A1(n_7182_o_0),
    .A2(net46),
    .B(net79),
    .C(n_7224_o_0),
    .Y(n_7620_o_0));
 AOI31xp33_ASAP7_75t_R n_7621 (.A1(n_7205_o_0),
    .A2(n_7220_o_0),
    .A3(net46),
    .B(n_7620_o_0),
    .Y(n_7621_o_0));
 OAI21xp33_ASAP7_75t_R n_7622 (.A1(n_7240_o_0),
    .A2(n_7621_o_0),
    .B(n_7261_o_0),
    .Y(n_7622_o_0));
 AOI21xp33_ASAP7_75t_R n_7623 (.A1(n_7229_o_0),
    .A2(n_7619_o_0),
    .B(n_7622_o_0),
    .Y(n_7623_o_0));
 AOI21xp33_ASAP7_75t_R n_7624 (.A1(n_7611_o_0),
    .A2(n_7616_o_0),
    .B(n_7623_o_0),
    .Y(n_7624_o_0));
 MAJIxp5_ASAP7_75t_R n_7625 (.A(n_7201_o_0),
    .B(n_7182_o_0),
    .C(net46),
    .Y(n_7625_o_0));
 OAI22xp33_ASAP7_75t_R n_7626 (.A1(n_7543_o_0),
    .A2(n_7482_o_0),
    .B1(n_7224_o_0),
    .B2(n_7625_o_0),
    .Y(n_7626_o_0));
 OAI21xp33_ASAP7_75t_R n_7627 (.A1(net46),
    .A2(n_7220_o_0),
    .B(n_7219_o_0),
    .Y(n_7627_o_0));
 AOI21xp33_ASAP7_75t_R n_7628 (.A1(net46),
    .A2(n_7182_o_0),
    .B(n_7627_o_0),
    .Y(n_7628_o_0));
 AOI211xp5_ASAP7_75t_R n_7629 (.A1(n_7224_o_0),
    .A2(n_7337_o_0),
    .B(n_7628_o_0),
    .C(n_7271_o_0),
    .Y(n_7629_o_0));
 AOI21xp33_ASAP7_75t_R n_7630 (.A1(n_7229_o_0),
    .A2(n_7626_o_0),
    .B(n_7629_o_0),
    .Y(n_7630_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7631 (.A1(n_7201_o_0),
    .A2(n_7224_o_0),
    .B(n_7339_o_0),
    .C(n_7353_o_0),
    .Y(n_7631_o_0));
 AOI21xp33_ASAP7_75t_R n_7632 (.A1(n_7240_o_0),
    .A2(n_7631_o_0),
    .B(n_7261_o_0),
    .Y(n_7632_o_0));
 OAI21xp33_ASAP7_75t_R n_7633 (.A1(n_7409_o_0),
    .A2(n_7336_o_0),
    .B(n_7219_o_0),
    .Y(n_7633_o_0));
 NAND3xp33_ASAP7_75t_R n_7634 (.A(n_7633_o_0),
    .B(n_7217_o_0),
    .C(n_7213_o_0),
    .Y(n_7634_o_0));
 AOI21xp33_ASAP7_75t_R n_7635 (.A1(n_7632_o_0),
    .A2(n_7634_o_0),
    .B(n_7367_o_0),
    .Y(n_7635_o_0));
 OAI21xp33_ASAP7_75t_R n_7636 (.A1(n_7279_o_0),
    .A2(n_7630_o_0),
    .B(n_7635_o_0),
    .Y(n_7636_o_0));
 OAI21xp33_ASAP7_75t_R n_7637 (.A1(n_7326_o_0),
    .A2(n_7624_o_0),
    .B(n_7636_o_0),
    .Y(n_7637_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7638 (.A1(n_7284_o_0),
    .A2(n_7249_o_0),
    .B(n_7255_o_0),
    .C(n_7241_o_0),
    .Y(n_7638_o_0));
 AOI21xp33_ASAP7_75t_R n_7639 (.A1(n_7229_o_0),
    .A2(n_7427_o_0),
    .B(n_7260_o_0),
    .Y(n_7639_o_0));
 OA21x2_ASAP7_75t_R n_7640 (.A1(n_7202_o_0),
    .A2(net46),
    .B(n_7382_o_0),
    .Y(n_7640_o_0));
 NAND2xp33_ASAP7_75t_R n_7641 (.A(n_7201_o_0),
    .B(n_7196_o_0),
    .Y(n_7641_o_0));
 OAI21xp33_ASAP7_75t_R n_7642 (.A1(n_7201_o_0),
    .A2(n_7196_o_0),
    .B(n_7641_o_0),
    .Y(n_7642_o_0));
 AO221x1_ASAP7_75t_R n_7643 (.A1(n_7151_o_0),
    .A2(n_7642_o_0),
    .B1(n_7205_o_0),
    .B2(n_7591_o_0),
    .C(n_7241_o_0),
    .Y(n_7643_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7644 (.A1(n_7331_o_0),
    .A2(n_7640_o_0),
    .B(n_7643_o_0),
    .C(n_7134_o_0),
    .Y(n_7644_o_0));
 AOI21xp33_ASAP7_75t_R n_7645 (.A1(n_7638_o_0),
    .A2(n_7639_o_0),
    .B(n_7644_o_0),
    .Y(n_7645_o_0));
 AOI21xp33_ASAP7_75t_R n_7646 (.A1(n_7450_o_0),
    .A2(n_7345_o_0),
    .B(n_7399_o_0),
    .Y(n_7646_o_0));
 OAI21xp33_ASAP7_75t_R n_7647 (.A1(n_7182_o_0),
    .A2(n_7224_o_0),
    .B(n_7201_o_0),
    .Y(n_7647_o_0));
 NAND3xp33_ASAP7_75t_R n_7648 (.A(n_7229_o_0),
    .B(n_7377_o_0),
    .C(n_7647_o_0),
    .Y(n_7648_o_0));
 OAI21xp33_ASAP7_75t_R n_7649 (.A1(n_7240_o_0),
    .A2(n_7646_o_0),
    .B(n_7648_o_0),
    .Y(n_7649_o_0));
 OAI211xp5_ASAP7_75t_R n_7650 (.A1(n_7436_o_0),
    .A2(n_7250_o_0),
    .B(n_7213_o_0),
    .C(n_7389_o_0),
    .Y(n_7650_o_0));
 OAI211xp5_ASAP7_75t_R n_7651 (.A1(n_7613_o_0),
    .A2(n_7151_o_0),
    .B(n_7570_o_0),
    .C(n_7229_o_0),
    .Y(n_7651_o_0));
 AOI31xp33_ASAP7_75t_R n_7652 (.A1(n_7261_o_0),
    .A2(n_7650_o_0),
    .A3(n_7651_o_0),
    .B(n_7327_o_0),
    .Y(n_7652_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7653 (.A1(n_7134_o_0),
    .A2(n_7649_o_0),
    .B(n_7652_o_0),
    .C(n_7274_o_0),
    .Y(n_7653_o_0));
 OAI21xp33_ASAP7_75t_R n_7654 (.A1(n_7366_o_0),
    .A2(n_7645_o_0),
    .B(n_7653_o_0),
    .Y(n_7654_o_0));
 OAI21xp33_ASAP7_75t_R n_7655 (.A1(n_7275_o_0),
    .A2(n_7637_o_0),
    .B(n_7654_o_0),
    .Y(n_7655_o_0));
 NOR2xp33_ASAP7_75t_R n_7656 (.A(n_7201_o_0),
    .B(n_7377_o_0),
    .Y(n_7656_o_0));
 OAI321xp33_ASAP7_75t_R n_7657 (.A1(n_7219_o_0),
    .A2(n_7656_o_0),
    .A3(n_7283_o_0),
    .B1(n_7450_o_0),
    .B2(n_7263_o_0),
    .C(n_7279_o_0),
    .Y(n_7657_o_0));
 OAI31xp33_ASAP7_75t_R n_7658 (.A1(n_7279_o_0),
    .A2(n_7356_o_0),
    .A3(n_7476_o_0),
    .B(n_7657_o_0),
    .Y(n_7658_o_0));
 OAI22xp33_ASAP7_75t_R n_7659 (.A1(n_7426_o_0),
    .A2(n_7224_o_0),
    .B1(n_7206_o_0),
    .B2(n_7656_o_0),
    .Y(n_7659_o_0));
 OAI21xp33_ASAP7_75t_R n_7660 (.A1(net23),
    .A2(n_7389_o_0),
    .B(n_7279_o_0),
    .Y(n_7660_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7661 (.A1(n_7182_o_0),
    .A2(n_7205_o_0),
    .B(n_7660_o_0),
    .C(n_7241_o_0),
    .Y(n_7661_o_0));
 AOI21xp33_ASAP7_75t_R n_7662 (.A1(n_7261_o_0),
    .A2(n_7659_o_0),
    .B(n_7661_o_0),
    .Y(n_7662_o_0));
 AOI21xp33_ASAP7_75t_R n_7663 (.A1(n_7229_o_0),
    .A2(n_7658_o_0),
    .B(n_7662_o_0),
    .Y(n_7663_o_0));
 AOI211xp5_ASAP7_75t_R n_7664 (.A1(n_7216_o_0),
    .A2(n_7196_o_0),
    .B(n_7291_o_0),
    .C(n_7281_o_0),
    .Y(n_7664_o_0));
 AO21x1_ASAP7_75t_R n_7665 (.A1(n_7300_o_0),
    .A2(n_7196_o_0),
    .B(n_7306_o_0),
    .Y(n_7665_o_0));
 OAI21xp33_ASAP7_75t_R n_7666 (.A1(n_7205_o_0),
    .A2(n_7664_o_0),
    .B(n_7665_o_0),
    .Y(n_7666_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7667 (.A1(n_7242_o_0),
    .A2(n_7402_o_0),
    .B(n_7392_o_0),
    .C(n_7260_o_0),
    .Y(n_7667_o_0));
 AOI21xp33_ASAP7_75t_R n_7668 (.A1(n_7279_o_0),
    .A2(n_7666_o_0),
    .B(n_7667_o_0),
    .Y(n_7668_o_0));
 NAND2xp33_ASAP7_75t_R n_7669 (.A(n_7543_o_0),
    .B(n_7536_o_0),
    .Y(n_7669_o_0));
 OA21x2_ASAP7_75t_R n_7670 (.A1(n_7543_o_0),
    .A2(n_7482_o_0),
    .B(n_7261_o_0),
    .Y(n_7670_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7671 (.A1(net23),
    .A2(n_7338_o_0),
    .B(n_7670_o_0),
    .C(n_7213_o_0),
    .Y(n_7671_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7672 (.A1(n_7134_o_0),
    .A2(n_7669_o_0),
    .B(n_7671_o_0),
    .C(n_7367_o_0),
    .Y(n_7672_o_0));
 OAI21xp33_ASAP7_75t_R n_7673 (.A1(n_7240_o_0),
    .A2(n_7668_o_0),
    .B(n_7672_o_0),
    .Y(n_7673_o_0));
 OAI21xp33_ASAP7_75t_R n_7674 (.A1(n_7366_o_0),
    .A2(n_7663_o_0),
    .B(n_7673_o_0),
    .Y(n_7674_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7675 (.A1(n_7224_o_0),
    .A2(n_7344_o_0),
    .B(n_7268_o_0),
    .C(n_7241_o_0),
    .Y(n_7675_o_0));
 AOI211xp5_ASAP7_75t_R n_7676 (.A1(n_7196_o_0),
    .A2(n_7179_o_0),
    .B(n_7151_o_0),
    .C(n_7201_o_0),
    .Y(n_7676_o_0));
 OAI211xp5_ASAP7_75t_R n_7677 (.A1(net46),
    .A2(n_7262_o_0),
    .B(n_7339_o_0),
    .C(n_7219_o_0),
    .Y(n_7677_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7678 (.A1(n_7219_o_0),
    .A2(n_7676_o_0),
    .B(n_7677_o_0),
    .C(n_7240_o_0),
    .Y(n_7678_o_0));
 OAI32xp33_ASAP7_75t_R n_7679 (.A1(n_7219_o_0),
    .A2(n_7409_o_0),
    .A3(n_7197_o_0),
    .B1(n_7224_o_0),
    .B2(n_7362_o_0),
    .Y(n_7679_o_0));
 AOI211xp5_ASAP7_75t_R n_7680 (.A1(n_7201_o_0),
    .A2(n_7196_o_0),
    .B(n_7281_o_0),
    .C(n_7219_o_0),
    .Y(n_7680_o_0));
 AOI31xp33_ASAP7_75t_R n_7681 (.A1(n_7151_o_0),
    .A2(n_7198_o_0),
    .A3(n_7613_o_0),
    .B(n_7680_o_0),
    .Y(n_7681_o_0));
 OAI321xp33_ASAP7_75t_R n_7682 (.A1(n_7679_o_0),
    .A2(n_7239_o_0),
    .A3(n_7564_o_0),
    .B1(n_7681_o_0),
    .B2(n_7240_o_0),
    .C(n_7261_o_0),
    .Y(n_7682_o_0));
 OAI31xp33_ASAP7_75t_R n_7683 (.A1(n_7261_o_0),
    .A2(n_7675_o_0),
    .A3(n_7678_o_0),
    .B(n_7682_o_0),
    .Y(n_7683_o_0));
 NAND2xp33_ASAP7_75t_R n_7684 (.A(n_7225_o_0),
    .B(n_7497_o_0),
    .Y(n_7684_o_0));
 OAI31xp33_ASAP7_75t_R n_7685 (.A1(n_7504_o_0),
    .A2(n_7291_o_0),
    .A3(n_7580_o_0),
    .B(n_7684_o_0),
    .Y(n_7685_o_0));
 OAI22xp33_ASAP7_75t_R n_7686 (.A1(n_7472_o_0),
    .A2(n_7482_o_0),
    .B1(n_7396_o_0),
    .B2(n_7373_o_0),
    .Y(n_7686_o_0));
 NOR3xp33_ASAP7_75t_R n_7687 (.A(n_7472_o_0),
    .B(n_7482_o_0),
    .C(n_7205_o_0),
    .Y(n_7687_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7688 (.A1(n_7205_o_0),
    .A2(n_7686_o_0),
    .B(n_7687_o_0),
    .C(n_7241_o_0),
    .D(n_7261_o_0),
    .Y(n_7688_o_0));
 OAI21xp33_ASAP7_75t_R n_7689 (.A1(n_7241_o_0),
    .A2(n_7685_o_0),
    .B(n_7688_o_0),
    .Y(n_7689_o_0));
 AOI22xp33_ASAP7_75t_R n_7690 (.A1(n_7339_o_0),
    .A2(n_7353_o_0),
    .B1(n_7205_o_0),
    .B2(n_7262_o_0),
    .Y(n_7690_o_0));
 OAI22xp33_ASAP7_75t_R n_7691 (.A1(n_7266_o_0),
    .A2(net46),
    .B1(n_7205_o_0),
    .B2(n_7506_o_0),
    .Y(n_7691_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7692 (.A1(n_7266_o_0),
    .A2(n_7267_o_0),
    .B(n_7691_o_0),
    .C(n_7240_o_0),
    .Y(n_7692_o_0));
 OAI211xp5_ASAP7_75t_R n_7693 (.A1(n_7229_o_0),
    .A2(n_7690_o_0),
    .B(n_7692_o_0),
    .C(n_7134_o_0),
    .Y(n_7693_o_0));
 AOI31xp33_ASAP7_75t_R n_7694 (.A1(n_7366_o_0),
    .A2(n_7689_o_0),
    .A3(n_7693_o_0),
    .B(n_7275_o_0),
    .Y(n_7694_o_0));
 OA21x2_ASAP7_75t_R n_7695 (.A1(n_7326_o_0),
    .A2(n_7683_o_0),
    .B(n_7694_o_0),
    .Y(n_7695_o_0));
 AOI21xp33_ASAP7_75t_R n_7696 (.A1(n_7519_o_0),
    .A2(n_7674_o_0),
    .B(n_7695_o_0),
    .Y(n_7696_o_0));
 INVx1_ASAP7_75t_R n_7697 (.A(_00642_),
    .Y(n_7697_o_0));
 XNOR2xp5_ASAP7_75t_R n_7698 (.A(_01082_),
    .B(_01121_),
    .Y(n_7698_o_0));
 XNOR2xp5_ASAP7_75t_R n_7699 (.A(n_7698_o_0),
    .B(n_3048_o_0),
    .Y(n_7699_o_0));
 NOR2xp33_ASAP7_75t_R n_7700 (.A(n_7697_o_0),
    .B(n_7699_o_0),
    .Y(n_7700_o_0));
 NOR2xp33_ASAP7_75t_R n_7701 (.A(_00659_),
    .B(net),
    .Y(n_7701_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7702 (.A1(n_7697_o_0),
    .A2(n_7699_o_0),
    .B(n_7700_o_0),
    .C(net),
    .D(n_7701_o_0),
    .Y(n_7702_o_0));
 XNOR2xp5_ASAP7_75t_R n_7703 (.A(_00875_),
    .B(n_7702_o_0),
    .Y(n_7703_o_0));
 XNOR2xp5_ASAP7_75t_R n_7704 (.A(_01121_),
    .B(n_3005_o_0),
    .Y(n_7704_o_0));
 NOR2xp33_ASAP7_75t_R n_7705 (.A(n_3011_o_0),
    .B(n_7704_o_0),
    .Y(n_7705_o_0));
 NOR2xp33_ASAP7_75t_R n_7706 (.A(_00660_),
    .B(net),
    .Y(n_7706_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7707 (.A1(n_3011_o_0),
    .A2(n_7704_o_0),
    .B(n_7705_o_0),
    .C(net),
    .D(n_7706_o_0),
    .Y(n_7707_o_0));
 XNOR2xp5_ASAP7_75t_R n_7708 (.A(_00874_),
    .B(n_7707_o_0),
    .Y(n_7708_o_0));
 NAND2xp33_ASAP7_75t_R n_7709 (.A(n_3113_o_0),
    .B(n_3135_o_0),
    .Y(n_7709_o_0));
 OAI21xp33_ASAP7_75t_R n_7710 (.A1(n_3113_o_0),
    .A2(n_3135_o_0),
    .B(n_7709_o_0),
    .Y(n_7710_o_0));
 NOR2xp33_ASAP7_75t_R n_7711 (.A(_01120_),
    .B(n_7710_o_0),
    .Y(n_7711_o_0));
 NOR2xp33_ASAP7_75t_R n_7712 (.A(_00661_),
    .B(net),
    .Y(n_7712_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7713 (.A1(n_7710_o_0),
    .A2(_01120_),
    .B(n_7711_o_0),
    .C(net),
    .D(n_7712_o_0),
    .Y(n_7713_o_0));
 XOR2xp5_ASAP7_75t_R n_7714 (.A(_00873_),
    .B(n_7713_o_0),
    .Y(n_7714_o_0));
 XNOR2xp5_ASAP7_75t_R n_7715 (.A(_01119_),
    .B(n_5516_o_0),
    .Y(n_7715_o_0));
 XNOR2xp5_ASAP7_75t_R n_7716 (.A(_00642_),
    .B(_01118_),
    .Y(n_7716_o_0));
 XNOR2xp5_ASAP7_75t_R n_7717 (.A(n_3004_o_0),
    .B(n_7716_o_0),
    .Y(n_7717_o_0));
 XNOR2xp5_ASAP7_75t_R n_7718 (.A(n_7715_o_0),
    .B(n_7717_o_0),
    .Y(n_7718_o_0));
 OR2x2_ASAP7_75t_R n_7719 (.A(_00662_),
    .B(net77),
    .Y(n_7719_o_0));
 OAI21xp33_ASAP7_75t_R n_7720 (.A1(net1),
    .A2(n_7718_o_0),
    .B(n_7719_o_0),
    .Y(n_7720_o_0));
 NAND2xp33_ASAP7_75t_R n_7721 (.A(_00872_),
    .B(n_7720_o_0),
    .Y(n_7721_o_0));
 OAI21xp5_ASAP7_75t_R n_7722 (.A1(_00872_),
    .A2(n_7720_o_0),
    .B(n_7721_o_0),
    .Y(n_7722_o_0));
 INVx1_ASAP7_75t_R n_7723 (.A(n_7722_o_0),
    .Y(n_7723_o_0));
 INVx1_ASAP7_75t_R n_7724 (.A(_00871_),
    .Y(n_7724_o_0));
 XNOR2xp5_ASAP7_75t_R n_7725 (.A(_00999_),
    .B(_01039_),
    .Y(n_7725_o_0));
 XOR2xp5_ASAP7_75t_R n_7726 (.A(_00642_),
    .B(_01117_),
    .Y(n_7726_o_0));
 XNOR2xp5_ASAP7_75t_R n_7727 (.A(n_7725_o_0),
    .B(n_7726_o_0),
    .Y(n_7727_o_0));
 XNOR2xp5_ASAP7_75t_R n_7728 (.A(_00643_),
    .B(_01078_),
    .Y(n_7728_o_0));
 XNOR2xp5_ASAP7_75t_R n_7729 (.A(_01118_),
    .B(n_7728_o_0),
    .Y(n_7729_o_0));
 NOR2xp33_ASAP7_75t_R n_7730 (.A(n_7729_o_0),
    .B(n_7727_o_0),
    .Y(n_7730_o_0));
 NOR2xp33_ASAP7_75t_R n_7731 (.A(_00663_),
    .B(_00858_),
    .Y(n_7731_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7732 (.A1(n_7727_o_0),
    .A2(n_7729_o_0),
    .B(n_7730_o_0),
    .C(net39),
    .D(n_7731_o_0),
    .Y(n_7732_o_0));
 NOR2xp33_ASAP7_75t_R n_7733 (.A(_01118_),
    .B(n_5491_o_0),
    .Y(n_7733_o_0));
 XNOR2xp5_ASAP7_75t_R n_7734 (.A(_00642_),
    .B(_01117_),
    .Y(n_7734_o_0));
 XNOR2xp5_ASAP7_75t_R n_7735 (.A(n_7725_o_0),
    .B(n_7734_o_0),
    .Y(n_7735_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7736 (.A1(_01118_),
    .A2(n_5491_o_0),
    .B(n_7733_o_0),
    .C(n_7735_o_0),
    .Y(n_7736_o_0));
 NAND2xp33_ASAP7_75t_R n_7737 (.A(n_7729_o_0),
    .B(n_7727_o_0),
    .Y(n_7737_o_0));
 INVx1_ASAP7_75t_R n_7738 (.A(n_7731_o_0),
    .Y(n_7738_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7739 (.A1(n_7736_o_0),
    .A2(n_7737_o_0),
    .B(net1),
    .C(n_7738_o_0),
    .D(n_7724_o_0),
    .Y(n_7739_o_0));
 AOI21xp5_ASAP7_75t_R n_7740 (.A1(n_7724_o_0),
    .A2(n_7732_o_0),
    .B(n_7739_o_0),
    .Y(n_7740_o_0));
 INVx1_ASAP7_75t_R n_7741 (.A(_00870_),
    .Y(n_7741_o_0));
 XNOR2xp5_ASAP7_75t_R n_7742 (.A(_00998_),
    .B(_01038_),
    .Y(n_7742_o_0));
 NAND2xp33_ASAP7_75t_R n_7743 (.A(_01117_),
    .B(n_7742_o_0),
    .Y(n_7743_o_0));
 OAI21xp33_ASAP7_75t_R n_7744 (.A1(_01117_),
    .A2(n_7742_o_0),
    .B(n_7743_o_0),
    .Y(n_7744_o_0));
 XOR2xp5_ASAP7_75t_R n_7745 (.A(_00998_),
    .B(_01038_),
    .Y(n_7745_o_0));
 INVx1_ASAP7_75t_R n_7746 (.A(_01117_),
    .Y(n_7746_o_0));
 NOR2xp33_ASAP7_75t_R n_7747 (.A(n_7746_o_0),
    .B(n_7745_o_0),
    .Y(n_7747_o_0));
 AOI211xp5_ASAP7_75t_R n_7748 (.A1(n_7745_o_0),
    .A2(n_7746_o_0),
    .B(n_7747_o_0),
    .C(n_5445_o_0),
    .Y(n_7748_o_0));
 NOR2xp33_ASAP7_75t_R n_7749 (.A(_00572_),
    .B(net77),
    .Y(n_7749_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7750 (.A1(n_5445_o_0),
    .A2(n_7744_o_0),
    .B(n_7748_o_0),
    .C(net39),
    .D(n_7749_o_0),
    .Y(n_7750_o_0));
 OAI211xp5_ASAP7_75t_R n_7751 (.A1(_01117_),
    .A2(n_7742_o_0),
    .B(n_7743_o_0),
    .C(n_5450_o_0),
    .Y(n_7751_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7752 (.A1(n_7745_o_0),
    .A2(n_7746_o_0),
    .B(n_7747_o_0),
    .C(n_5445_o_0),
    .Y(n_7752_o_0));
 INVx1_ASAP7_75t_R n_7753 (.A(n_7749_o_0),
    .Y(n_7753_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7754 (.A1(n_7751_o_0),
    .A2(n_7752_o_0),
    .B(net3),
    .C(n_7753_o_0),
    .D(n_7741_o_0),
    .Y(n_7754_o_0));
 AO21x2_ASAP7_75t_R n_7755 (.A1(n_7741_o_0),
    .A2(n_7750_o_0),
    .B(n_7754_o_0),
    .Y(n_7755_o_0));
 XNOR2xp5_ASAP7_75t_R n_7756 (.A(_00996_),
    .B(_01036_),
    .Y(n_7756_o_0));
 INVx1_ASAP7_75t_R n_7757 (.A(_00643_),
    .Y(n_7757_o_0));
 NOR2xp33_ASAP7_75t_R n_7758 (.A(n_7757_o_0),
    .B(n_7756_o_0),
    .Y(n_7758_o_0));
 XNOR2xp5_ASAP7_75t_R n_7759 (.A(_00642_),
    .B(_01115_),
    .Y(n_7759_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7760 (.A1(n_7756_o_0),
    .A2(n_7757_o_0),
    .B(n_7758_o_0),
    .C(n_7759_o_0),
    .Y(n_7760_o_0));
 NAND2xp33_ASAP7_75t_R n_7761 (.A(n_7757_o_0),
    .B(n_7756_o_0),
    .Y(n_7761_o_0));
 XOR2xp5_ASAP7_75t_R n_7762 (.A(_00642_),
    .B(_01115_),
    .Y(n_7762_o_0));
 OAI211xp5_ASAP7_75t_R n_7763 (.A1(n_7756_o_0),
    .A2(n_7757_o_0),
    .B(n_7761_o_0),
    .C(n_7762_o_0),
    .Y(n_7763_o_0));
 OR2x2_ASAP7_75t_R n_7764 (.A(_00570_),
    .B(net39),
    .Y(n_7764_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7765 (.A1(n_7760_o_0),
    .A2(n_7763_o_0),
    .B(net5),
    .C(n_7764_o_0),
    .Y(n_7765_o_0));
 INVx1_ASAP7_75t_R n_7766 (.A(n_7765_o_0),
    .Y(n_7766_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7767 (.A1(n_7763_o_0),
    .A2(n_7760_o_0),
    .B(net5),
    .C(n_7764_o_0),
    .D(_00868_),
    .Y(n_7767_o_0));
 AOI21x1_ASAP7_75t_R n_7768 (.A1(_00868_),
    .A2(n_7766_o_0),
    .B(n_7767_o_0),
    .Y(n_7768_o_0));
 NAND2xp33_ASAP7_75t_R n_7769 (.A(n_3035_o_0),
    .B(n_5444_o_0),
    .Y(n_7769_o_0));
 XNOR2xp5_ASAP7_75t_R n_7770 (.A(_01116_),
    .B(n_7759_o_0),
    .Y(n_7770_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7771 (.A1(n_5444_o_0),
    .A2(n_3035_o_0),
    .B(n_7769_o_0),
    .C(n_7770_o_0),
    .Y(n_7771_o_0));
 XNOR2xp5_ASAP7_75t_R n_7772 (.A(n_3067_o_0),
    .B(n_7759_o_0),
    .Y(n_7772_o_0));
 OAI21xp33_ASAP7_75t_R n_7773 (.A1(n_5444_o_0),
    .A2(n_3035_o_0),
    .B(n_7769_o_0),
    .Y(n_7773_o_0));
 OAI21xp33_ASAP7_75t_R n_7774 (.A1(n_7772_o_0),
    .A2(n_7773_o_0),
    .B(_00858_),
    .Y(n_7774_o_0));
 NOR2xp33_ASAP7_75t_R n_7775 (.A(n_7771_o_0),
    .B(n_7774_o_0),
    .Y(n_7775_o_0));
 INVx1_ASAP7_75t_R n_7776 (.A(_00569_),
    .Y(n_7776_o_0));
 INVx1_ASAP7_75t_R n_7777 (.A(_00869_),
    .Y(n_7777_o_0));
 OA221x2_ASAP7_75t_R n_7778 (.A1(net),
    .A2(n_7776_o_0),
    .B1(n_7774_o_0),
    .B2(n_7771_o_0),
    .C(n_7777_o_0),
    .Y(n_7778_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_7779 (.A1(net9),
    .A2(_00569_),
    .B(n_7775_o_0),
    .C(_00869_),
    .D(n_7778_o_0),
    .Y(n_7779_o_0));
 NOR2xp33_ASAP7_75t_R n_7780 (.A(n_7768_o_0),
    .B(n_7779_o_0),
    .Y(n_7780_o_0));
 NOR2xp33_ASAP7_75t_R n_7781 (.A(n_7755_o_0),
    .B(n_7780_o_0),
    .Y(n_7781_o_0));
 AO21x1_ASAP7_75t_R n_7782 (.A1(n_7766_o_0),
    .A2(_00868_),
    .B(n_7767_o_0),
    .Y(n_7782_o_0));
 NAND2xp33_ASAP7_75t_R n_7783 (.A(n_7779_o_0),
    .B(n_7782_o_0),
    .Y(n_7783_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7784 (.A1(n_7737_o_0),
    .A2(n_7736_o_0),
    .B(net5),
    .C(n_7738_o_0),
    .Y(n_7784_o_0));
 NAND2xp33_ASAP7_75t_R n_7785 (.A(n_7724_o_0),
    .B(n_7784_o_0),
    .Y(n_7785_o_0));
 OAI21xp5_ASAP7_75t_R n_7786 (.A1(n_7724_o_0),
    .A2(n_7784_o_0),
    .B(n_7785_o_0),
    .Y(n_7786_o_0));
 NOR2xp33_ASAP7_75t_R n_7787 (.A(n_3035_o_0),
    .B(n_5444_o_0),
    .Y(n_7787_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7788 (.A1(n_5444_o_0),
    .A2(n_3035_o_0),
    .B(n_7787_o_0),
    .C(n_7772_o_0),
    .Y(n_7788_o_0));
 OAI211xp5_ASAP7_75t_R n_7789 (.A1(n_7772_o_0),
    .A2(n_7773_o_0),
    .B(n_7788_o_0),
    .C(net39),
    .Y(n_7789_o_0));
 NAND2xp33_ASAP7_75t_R n_7790 (.A(_00569_),
    .B(net5),
    .Y(n_7790_o_0));
 OAI221xp5_ASAP7_75t_R n_7791 (.A1(net39),
    .A2(n_7776_o_0),
    .B1(n_7771_o_0),
    .B2(n_7774_o_0),
    .C(n_7777_o_0),
    .Y(n_7791_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7792 (.A1(n_7789_o_0),
    .A2(n_7790_o_0),
    .B(n_7777_o_0),
    .C(n_7791_o_0),
    .Y(n_7792_o_0));
 NAND4xp25_ASAP7_75t_R n_7793 (.A(n_7782_o_0),
    .B(n_7740_o_0),
    .C(n_7755_o_0),
    .D(net34),
    .Y(n_7793_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7794 (.A1(n_7783_o_0),
    .A2(n_7755_o_0),
    .B(n_7786_o_0),
    .C(n_7793_o_0),
    .Y(n_7794_o_0));
 AO21x1_ASAP7_75t_R n_7795 (.A1(n_7740_o_0),
    .A2(n_7781_o_0),
    .B(n_7794_o_0),
    .Y(n_7795_o_0));
 AOI21x1_ASAP7_75t_R n_7796 (.A1(n_7741_o_0),
    .A2(n_7750_o_0),
    .B(n_7754_o_0),
    .Y(n_7796_o_0));
 NOR2xp33_ASAP7_75t_R n_7797 (.A(n_7796_o_0),
    .B(n_7768_o_0),
    .Y(n_7797_o_0));
 NAND2xp33_ASAP7_75t_R n_7798 (.A(n_7792_o_0),
    .B(n_7768_o_0),
    .Y(n_7798_o_0));
 NOR2xp33_ASAP7_75t_R n_7799 (.A(n_7755_o_0),
    .B(n_7798_o_0),
    .Y(n_7799_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7800 (.A1(_00868_),
    .A2(n_7766_o_0),
    .B(n_7767_o_0),
    .C(n_7792_o_0),
    .Y(n_7800_o_0));
 OAI21xp33_ASAP7_75t_R n_7801 (.A1(n_7782_o_0),
    .A2(n_7792_o_0),
    .B(n_7800_o_0),
    .Y(n_7801_o_0));
 OAI21xp33_ASAP7_75t_R n_7802 (.A1(n_7796_o_0),
    .A2(net97),
    .B(n_7786_o_0),
    .Y(n_7802_o_0));
 INVx1_ASAP7_75t_R n_7803 (.A(n_7802_o_0),
    .Y(n_7803_o_0));
 OAI21xp33_ASAP7_75t_R n_7804 (.A1(n_7755_o_0),
    .A2(n_7801_o_0),
    .B(n_7803_o_0),
    .Y(n_7804_o_0));
 OAI311xp33_ASAP7_75t_R n_7805 (.A1(n_7740_o_0),
    .A2(n_7797_o_0),
    .A3(n_7799_o_0),
    .B1(n_7723_o_0),
    .C1(n_7804_o_0),
    .Y(n_7805_o_0));
 OAI21xp33_ASAP7_75t_R n_7806 (.A1(n_7723_o_0),
    .A2(n_7795_o_0),
    .B(n_7805_o_0),
    .Y(n_7806_o_0));
 NAND2xp33_ASAP7_75t_R n_7807 (.A(n_7755_o_0),
    .B(n_7740_o_0),
    .Y(n_7807_o_0));
 NAND2xp33_ASAP7_75t_R n_7808 (.A(n_7768_o_0),
    .B(n_7779_o_0),
    .Y(n_7808_o_0));
 XNOR2xp5_ASAP7_75t_R n_7809 (.A(_00871_),
    .B(n_7784_o_0),
    .Y(n_7809_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7810 (.A1(n_7808_o_0),
    .A2(n_7800_o_0),
    .B(n_7796_o_0),
    .C(n_7809_o_0),
    .Y(n_7810_o_0));
 OAI211xp5_ASAP7_75t_R n_7811 (.A1(n_7807_o_0),
    .A2(n_7798_o_0),
    .B(n_7810_o_0),
    .C(n_7722_o_0),
    .Y(n_7811_o_0));
 NAND2xp5_ASAP7_75t_R n_7812 (.A(n_7779_o_0),
    .B(n_7768_o_0),
    .Y(n_7812_o_0));
 NOR2xp33_ASAP7_75t_R n_7813 (.A(n_7755_o_0),
    .B(n_7768_o_0),
    .Y(n_7813_o_0));
 INVx1_ASAP7_75t_R n_7814 (.A(n_7813_o_0),
    .Y(n_7814_o_0));
 AO21x1_ASAP7_75t_R n_7815 (.A1(n_5491_o_0),
    .A2(_01118_),
    .B(n_7733_o_0),
    .Y(n_7815_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7816 (.A1(n_7735_o_0),
    .A2(n_7815_o_0),
    .B(n_7736_o_0),
    .C(net2),
    .Y(n_7816_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7817 (.A1(net2),
    .A2(n_7731_o_0),
    .B(n_7816_o_0),
    .C(_00871_),
    .Y(n_7817_o_0));
 OAI21xp5_ASAP7_75t_R n_7818 (.A1(_00871_),
    .A2(n_7784_o_0),
    .B(n_7817_o_0),
    .Y(n_7818_o_0));
 OAI211xp5_ASAP7_75t_R n_7819 (.A1(n_7812_o_0),
    .A2(n_7796_o_0),
    .B(n_7814_o_0),
    .C(n_7818_o_0),
    .Y(n_7819_o_0));
 NAND2xp33_ASAP7_75t_R n_7820 (.A(n_7723_o_0),
    .B(n_7819_o_0),
    .Y(n_7820_o_0));
 OAI211xp5_ASAP7_75t_R n_7821 (.A1(_00871_),
    .A2(n_7784_o_0),
    .B(n_7817_o_0),
    .C(n_7796_o_0),
    .Y(n_7821_o_0));
 XOR2xp5_ASAP7_75t_R n_7822 (.A(_00873_),
    .B(n_7713_o_0),
    .Y(n_7822_o_0));
 INVx1_ASAP7_75t_R n_7823 (.A(n_7822_o_0),
    .Y(n_7823_o_0));
 OAI21xp33_ASAP7_75t_R n_7824 (.A1(n_7783_o_0),
    .A2(n_7821_o_0),
    .B(n_7823_o_0),
    .Y(n_7824_o_0));
 AOI21xp33_ASAP7_75t_R n_7825 (.A1(n_7811_o_0),
    .A2(n_7820_o_0),
    .B(n_7824_o_0),
    .Y(n_7825_o_0));
 AOI21xp33_ASAP7_75t_R n_7826 (.A1(n_7714_o_0),
    .A2(n_7806_o_0),
    .B(n_7825_o_0),
    .Y(n_7826_o_0));
 NOR2xp33_ASAP7_75t_R n_7827 (.A(n_7792_o_0),
    .B(n_7768_o_0),
    .Y(n_7827_o_0));
 NOR2xp33_ASAP7_75t_R n_7828 (.A(n_7827_o_0),
    .B(n_7807_o_0),
    .Y(n_7828_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7829 (.A1(net2),
    .A2(_00569_),
    .B(n_7775_o_0),
    .C(_00869_),
    .Y(n_7829_o_0));
 AOI21xp33_ASAP7_75t_R n_7830 (.A1(n_7791_o_0),
    .A2(n_7829_o_0),
    .B(n_7782_o_0),
    .Y(n_7830_o_0));
 NOR2xp33_ASAP7_75t_R n_7831 (.A(n_7821_o_0),
    .B(n_7830_o_0),
    .Y(n_7831_o_0));
 NAND2xp33_ASAP7_75t_R n_7832 (.A(n_7792_o_0),
    .B(n_7782_o_0),
    .Y(n_7832_o_0));
 OAI31xp33_ASAP7_75t_R n_7833 (.A1(n_7796_o_0),
    .A2(n_7832_o_0),
    .A3(n_7786_o_0),
    .B(n_7722_o_0),
    .Y(n_7833_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7834 (.A1(n_7768_o_0),
    .A2(net97),
    .B(n_7755_o_0),
    .C(n_7809_o_0),
    .Y(n_7834_o_0));
 INVx1_ASAP7_75t_R n_7835 (.A(_00872_),
    .Y(n_7835_o_0));
 NAND2xp33_ASAP7_75t_R n_7836 (.A(n_7835_o_0),
    .B(n_7720_o_0),
    .Y(n_7836_o_0));
 OAI21xp5_ASAP7_75t_R n_7837 (.A1(n_7835_o_0),
    .A2(n_7720_o_0),
    .B(n_7836_o_0),
    .Y(n_7837_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7838 (.A1(n_7755_o_0),
    .A2(n_7827_o_0),
    .B(n_7834_o_0),
    .C(n_7837_o_0),
    .Y(n_7838_o_0));
 INVx1_ASAP7_75t_R n_7839 (.A(n_7838_o_0),
    .Y(n_7839_o_0));
 OAI21xp33_ASAP7_75t_R n_7840 (.A1(n_7832_o_0),
    .A2(n_7807_o_0),
    .B(n_7839_o_0),
    .Y(n_7840_o_0));
 OAI31xp33_ASAP7_75t_R n_7841 (.A1(n_7828_o_0),
    .A2(n_7831_o_0),
    .A3(n_7833_o_0),
    .B(n_7840_o_0),
    .Y(n_7841_o_0));
 AOI21xp33_ASAP7_75t_R n_7842 (.A1(n_7791_o_0),
    .A2(n_7829_o_0),
    .B(n_7768_o_0),
    .Y(n_7842_o_0));
 AOI211xp5_ASAP7_75t_R n_7843 (.A1(n_7768_o_0),
    .A2(n_7779_o_0),
    .B(n_7842_o_0),
    .C(n_7755_o_0),
    .Y(n_7843_o_0));
 OAI21xp33_ASAP7_75t_R n_7844 (.A1(n_7796_o_0),
    .A2(net34),
    .B(n_7818_o_0),
    .Y(n_7844_o_0));
 OAI21xp33_ASAP7_75t_R n_7845 (.A1(n_7809_o_0),
    .A2(n_7843_o_0),
    .B(n_7844_o_0),
    .Y(n_7845_o_0));
 AOI21xp33_ASAP7_75t_R n_7846 (.A1(n_7722_o_0),
    .A2(n_7845_o_0),
    .B(n_7714_o_0),
    .Y(n_7846_o_0));
 OAI321xp33_ASAP7_75t_R n_7847 (.A1(net34),
    .A2(n_7821_o_0),
    .A3(n_7768_o_0),
    .B1(n_7807_o_0),
    .B2(n_7827_o_0),
    .C(n_7837_o_0),
    .Y(n_7847_o_0));
 INVx1_ASAP7_75t_R n_7848 (.A(n_7847_o_0),
    .Y(n_7848_o_0));
 AOI21xp33_ASAP7_75t_R n_7849 (.A1(n_7792_o_0),
    .A2(n_7782_o_0),
    .B(n_7796_o_0),
    .Y(n_7849_o_0));
 NAND2xp33_ASAP7_75t_R n_7850 (.A(n_7796_o_0),
    .B(n_7768_o_0),
    .Y(n_7850_o_0));
 INVx1_ASAP7_75t_R n_7851 (.A(n_7850_o_0),
    .Y(n_7851_o_0));
 OAI21xp33_ASAP7_75t_R n_7852 (.A1(n_7849_o_0),
    .A2(n_7851_o_0),
    .B(n_7809_o_0),
    .Y(n_7852_o_0));
 OAI211xp5_ASAP7_75t_R n_7853 (.A1(n_7832_o_0),
    .A2(n_7821_o_0),
    .B(n_7848_o_0),
    .C(n_7852_o_0),
    .Y(n_7853_o_0));
 NAND2xp33_ASAP7_75t_R n_7854 (.A(_00874_),
    .B(n_7707_o_0),
    .Y(n_7854_o_0));
 OAI21xp33_ASAP7_75t_R n_7855 (.A1(_00874_),
    .A2(n_7707_o_0),
    .B(n_7854_o_0),
    .Y(n_7855_o_0));
 INVx1_ASAP7_75t_R n_7856 (.A(n_7855_o_0),
    .Y(n_7856_o_0));
 AOI21xp33_ASAP7_75t_R n_7857 (.A1(n_7846_o_0),
    .A2(n_7853_o_0),
    .B(n_7856_o_0),
    .Y(n_7857_o_0));
 OAI21xp33_ASAP7_75t_R n_7858 (.A1(n_7823_o_0),
    .A2(n_7841_o_0),
    .B(n_7857_o_0),
    .Y(n_7858_o_0));
 OAI21xp33_ASAP7_75t_R n_7859 (.A1(n_7708_o_0),
    .A2(n_7826_o_0),
    .B(n_7858_o_0),
    .Y(n_7859_o_0));
 INVx1_ASAP7_75t_R n_7860 (.A(n_7708_o_0),
    .Y(n_7860_o_0));
 NOR2xp33_ASAP7_75t_R n_7861 (.A(n_7768_o_0),
    .B(n_7779_o_0),
    .Y(n_7861_o_0));
 INVx1_ASAP7_75t_R n_7862 (.A(n_7861_o_0),
    .Y(n_7862_o_0));
 OAI21xp33_ASAP7_75t_R n_7863 (.A1(n_7796_o_0),
    .A2(n_7782_o_0),
    .B(n_7786_o_0),
    .Y(n_7863_o_0));
 INVx1_ASAP7_75t_R n_7864 (.A(n_7863_o_0),
    .Y(n_7864_o_0));
 NAND2xp33_ASAP7_75t_R n_7865 (.A(n_7755_o_0),
    .B(n_7768_o_0),
    .Y(n_7865_o_0));
 INVx1_ASAP7_75t_R n_7866 (.A(n_7865_o_0),
    .Y(n_7866_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7867 (.A1(n_7861_o_0),
    .A2(n_7866_o_0),
    .B(n_7809_o_0),
    .C(n_7723_o_0),
    .Y(n_7867_o_0));
 INVx1_ASAP7_75t_R n_7868 (.A(n_7867_o_0),
    .Y(n_7868_o_0));
 OAI21xp33_ASAP7_75t_R n_7869 (.A1(n_7796_o_0),
    .A2(n_7798_o_0),
    .B(n_7809_o_0),
    .Y(n_7869_o_0));
 NOR2xp33_ASAP7_75t_R n_7870 (.A(n_7755_o_0),
    .B(n_7832_o_0),
    .Y(n_7870_o_0));
 NOR2xp33_ASAP7_75t_R n_7871 (.A(n_7755_o_0),
    .B(n_7812_o_0),
    .Y(n_7871_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7872 (.A1(n_7808_o_0),
    .A2(n_7800_o_0),
    .B(n_7796_o_0),
    .C(n_7740_o_0),
    .Y(n_7872_o_0));
 OAI221xp5_ASAP7_75t_R n_7873 (.A1(n_7869_o_0),
    .A2(n_7870_o_0),
    .B1(n_7871_o_0),
    .B2(n_7872_o_0),
    .C(n_7837_o_0),
    .Y(n_7873_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7874 (.A1(n_7862_o_0),
    .A2(n_7864_o_0),
    .B(n_7868_o_0),
    .C(n_7873_o_0),
    .Y(n_7874_o_0));
 INVx1_ASAP7_75t_R n_7875 (.A(n_7831_o_0),
    .Y(n_7875_o_0));
 NAND2xp33_ASAP7_75t_R n_7876 (.A(n_7740_o_0),
    .B(n_7849_o_0),
    .Y(n_7876_o_0));
 OAI211xp5_ASAP7_75t_R n_7877 (.A1(n_7810_o_0),
    .A2(n_7870_o_0),
    .B(n_7875_o_0),
    .C(n_7876_o_0),
    .Y(n_7877_o_0));
 AOI21xp33_ASAP7_75t_R n_7878 (.A1(n_7723_o_0),
    .A2(n_7877_o_0),
    .B(n_7822_o_0),
    .Y(n_7878_o_0));
 AOI22xp33_ASAP7_75t_R n_7879 (.A1(n_7808_o_0),
    .A2(n_7800_o_0),
    .B1(n_7755_o_0),
    .B2(n_7809_o_0),
    .Y(n_7879_o_0));
 NOR2xp33_ASAP7_75t_R n_7880 (.A(n_7809_o_0),
    .B(n_7801_o_0),
    .Y(n_7880_o_0));
 AOI31xp33_ASAP7_75t_R n_7881 (.A1(n_7755_o_0),
    .A2(n_7801_o_0),
    .A3(n_7786_o_0),
    .B(n_7837_o_0),
    .Y(n_7881_o_0));
 OAI221xp5_ASAP7_75t_R n_7882 (.A1(net96),
    .A2(n_7821_o_0),
    .B1(n_7879_o_0),
    .B2(n_7880_o_0),
    .C(n_7881_o_0),
    .Y(n_7882_o_0));
 AOI22xp33_ASAP7_75t_R n_7883 (.A1(n_7874_o_0),
    .A2(n_7714_o_0),
    .B1(n_7878_o_0),
    .B2(n_7882_o_0),
    .Y(n_7883_o_0));
 NOR3xp33_ASAP7_75t_R n_7884 (.A(n_7768_o_0),
    .B(net97),
    .C(n_7755_o_0),
    .Y(n_7884_o_0));
 INVx1_ASAP7_75t_R n_7885 (.A(n_7884_o_0),
    .Y(n_7885_o_0));
 AOI21xp33_ASAP7_75t_R n_7886 (.A1(n_7755_o_0),
    .A2(n_7783_o_0),
    .B(n_7786_o_0),
    .Y(n_7886_o_0));
 AOI21xp33_ASAP7_75t_R n_7887 (.A1(n_7885_o_0),
    .A2(n_7886_o_0),
    .B(n_7722_o_0),
    .Y(n_7887_o_0));
 OAI21xp33_ASAP7_75t_R n_7888 (.A1(n_7809_o_0),
    .A2(n_7813_o_0),
    .B(n_7887_o_0),
    .Y(n_7888_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7889 (.A1(n_7808_o_0),
    .A2(n_7800_o_0),
    .B(n_7796_o_0),
    .C(n_7809_o_0),
    .Y(n_7889_o_0));
 NOR2xp33_ASAP7_75t_R n_7890 (.A(n_7792_o_0),
    .B(n_7782_o_0),
    .Y(n_7890_o_0));
 NOR2xp33_ASAP7_75t_R n_7891 (.A(n_7755_o_0),
    .B(n_7890_o_0),
    .Y(n_7891_o_0));
 INVx1_ASAP7_75t_R n_7892 (.A(n_7797_o_0),
    .Y(n_7892_o_0));
 AOI21xp33_ASAP7_75t_R n_7893 (.A1(n_7796_o_0),
    .A2(n_7827_o_0),
    .B(n_7809_o_0),
    .Y(n_7893_o_0));
 AOI21xp33_ASAP7_75t_R n_7894 (.A1(n_7892_o_0),
    .A2(n_7893_o_0),
    .B(n_7837_o_0),
    .Y(n_7894_o_0));
 OAI21xp33_ASAP7_75t_R n_7895 (.A1(n_7889_o_0),
    .A2(n_7891_o_0),
    .B(n_7894_o_0),
    .Y(n_7895_o_0));
 NAND3xp33_ASAP7_75t_R n_7896 (.A(n_7888_o_0),
    .B(n_7895_o_0),
    .C(n_7714_o_0),
    .Y(n_7896_o_0));
 AOI21xp33_ASAP7_75t_R n_7897 (.A1(n_7768_o_0),
    .A2(n_7779_o_0),
    .B(n_7796_o_0),
    .Y(n_7897_o_0));
 NAND2xp33_ASAP7_75t_R n_7898 (.A(n_7755_o_0),
    .B(n_7792_o_0),
    .Y(n_7898_o_0));
 NAND2xp33_ASAP7_75t_R n_7899 (.A(n_7898_o_0),
    .B(n_7893_o_0),
    .Y(n_7899_o_0));
 OAI31xp33_ASAP7_75t_R n_7900 (.A1(n_7740_o_0),
    .A2(n_7813_o_0),
    .A3(n_7897_o_0),
    .B(n_7899_o_0),
    .Y(n_7900_o_0));
 OAI211xp5_ASAP7_75t_R n_7901 (.A1(n_7782_o_0),
    .A2(n_7796_o_0),
    .B(net34),
    .C(n_7740_o_0),
    .Y(n_7901_o_0));
 AOI31xp33_ASAP7_75t_R n_7902 (.A1(n_7723_o_0),
    .A2(n_7819_o_0),
    .A3(n_7901_o_0),
    .B(n_7822_o_0),
    .Y(n_7902_o_0));
 OAI21xp33_ASAP7_75t_R n_7903 (.A1(n_7837_o_0),
    .A2(n_7900_o_0),
    .B(n_7902_o_0),
    .Y(n_7903_o_0));
 NAND2xp33_ASAP7_75t_R n_7904 (.A(_00875_),
    .B(n_7702_o_0),
    .Y(n_7904_o_0));
 OAI21xp33_ASAP7_75t_R n_7905 (.A1(_00875_),
    .A2(n_7702_o_0),
    .B(n_7904_o_0),
    .Y(n_7905_o_0));
 INVx1_ASAP7_75t_R n_7906 (.A(n_7905_o_0),
    .Y(n_7906_o_0));
 AOI31xp33_ASAP7_75t_R n_7907 (.A1(n_7856_o_0),
    .A2(n_7896_o_0),
    .A3(n_7903_o_0),
    .B(n_7906_o_0),
    .Y(n_7907_o_0));
 OAI21xp33_ASAP7_75t_R n_7908 (.A1(n_7860_o_0),
    .A2(n_7883_o_0),
    .B(n_7907_o_0),
    .Y(n_7908_o_0));
 OAI21xp33_ASAP7_75t_R n_7909 (.A1(n_7703_o_0),
    .A2(n_7859_o_0),
    .B(n_7908_o_0),
    .Y(n_7909_o_0));
 INVx1_ASAP7_75t_R n_7910 (.A(n_7714_o_0),
    .Y(n_7910_o_0));
 NOR2xp33_ASAP7_75t_R n_7911 (.A(n_7755_o_0),
    .B(n_7740_o_0),
    .Y(n_7911_o_0));
 OAI21xp33_ASAP7_75t_R n_7912 (.A1(n_7802_o_0),
    .A2(n_7861_o_0),
    .B(n_7723_o_0),
    .Y(n_7912_o_0));
 AOI21xp33_ASAP7_75t_R n_7913 (.A1(n_7911_o_0),
    .A2(n_7783_o_0),
    .B(n_7912_o_0),
    .Y(n_7913_o_0));
 INVx1_ASAP7_75t_R n_7914 (.A(n_7889_o_0),
    .Y(n_7914_o_0));
 NAND2xp33_ASAP7_75t_R n_7915 (.A(n_7786_o_0),
    .B(n_7850_o_0),
    .Y(n_7915_o_0));
 INVx1_ASAP7_75t_R n_7916 (.A(n_7837_o_0),
    .Y(n_7916_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_7917 (.A1(n_7755_o_0),
    .A2(n_7783_o_0),
    .B(n_7915_o_0),
    .C(n_7916_o_0),
    .Y(n_7917_o_0));
 AOI21xp33_ASAP7_75t_R n_7918 (.A1(n_7814_o_0),
    .A2(n_7914_o_0),
    .B(n_7917_o_0),
    .Y(n_7918_o_0));
 AOI211xp5_ASAP7_75t_R n_7919 (.A1(n_7755_o_0),
    .A2(n_7812_o_0),
    .B(n_7880_o_0),
    .C(n_7879_o_0),
    .Y(n_7919_o_0));
 NOR2xp33_ASAP7_75t_R n_7920 (.A(n_7755_o_0),
    .B(net97),
    .Y(n_7920_o_0));
 AOI21xp33_ASAP7_75t_R n_7921 (.A1(n_7779_o_0),
    .A2(n_7782_o_0),
    .B(n_7755_o_0),
    .Y(n_7921_o_0));
 INVx1_ASAP7_75t_R n_7922 (.A(n_7921_o_0),
    .Y(n_7922_o_0));
 AOI21xp33_ASAP7_75t_R n_7923 (.A1(n_7922_o_0),
    .A2(n_7803_o_0),
    .B(n_7837_o_0),
    .Y(n_7923_o_0));
 OAI21xp33_ASAP7_75t_R n_7924 (.A1(n_7740_o_0),
    .A2(n_7920_o_0),
    .B(n_7923_o_0),
    .Y(n_7924_o_0));
 OAI211xp5_ASAP7_75t_R n_7925 (.A1(n_7919_o_0),
    .A2(n_7847_o_0),
    .B(n_7924_o_0),
    .C(n_7910_o_0),
    .Y(n_7925_o_0));
 OAI31xp33_ASAP7_75t_R n_7926 (.A1(n_7910_o_0),
    .A2(n_7913_o_0),
    .A3(n_7918_o_0),
    .B(n_7925_o_0),
    .Y(n_7926_o_0));
 NAND2xp33_ASAP7_75t_R n_7927 (.A(n_7768_o_0),
    .B(n_7779_o_0),
    .Y(n_7927_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7928 (.A1(n_7782_o_0),
    .A2(net34),
    .B(n_7800_o_0),
    .C(n_7755_o_0),
    .Y(n_7928_o_0));
 NOR2xp33_ASAP7_75t_R n_7929 (.A(n_7863_o_0),
    .B(n_7928_o_0),
    .Y(n_7929_o_0));
 AOI31xp33_ASAP7_75t_R n_7930 (.A1(n_7818_o_0),
    .A2(n_7892_o_0),
    .A3(n_7927_o_0),
    .B(n_7929_o_0),
    .Y(n_7930_o_0));
 OAI21xp33_ASAP7_75t_R n_7931 (.A1(n_7849_o_0),
    .A2(n_7915_o_0),
    .B(n_7916_o_0),
    .Y(n_7931_o_0));
 AOI21xp33_ASAP7_75t_R n_7932 (.A1(n_7885_o_0),
    .A2(n_7914_o_0),
    .B(n_7931_o_0),
    .Y(n_7932_o_0));
 AOI21xp33_ASAP7_75t_R n_7933 (.A1(n_7723_o_0),
    .A2(n_7930_o_0),
    .B(n_7932_o_0),
    .Y(n_7933_o_0));
 OAI211xp5_ASAP7_75t_R n_7934 (.A1(n_7782_o_0),
    .A2(n_7792_o_0),
    .B(n_7800_o_0),
    .C(n_7755_o_0),
    .Y(n_7934_o_0));
 OAI211xp5_ASAP7_75t_R n_7935 (.A1(n_7755_o_0),
    .A2(n_7812_o_0),
    .B(n_7934_o_0),
    .C(n_7818_o_0),
    .Y(n_7935_o_0));
 OAI31xp33_ASAP7_75t_R n_7936 (.A1(n_7796_o_0),
    .A2(n_7809_o_0),
    .A3(n_7783_o_0),
    .B(n_7935_o_0),
    .Y(n_7936_o_0));
 NAND4xp25_ASAP7_75t_R n_7937 (.A(n_7812_o_0),
    .B(n_7786_o_0),
    .C(n_7755_o_0),
    .D(n_7740_o_0),
    .Y(n_7937_o_0));
 NAND2xp33_ASAP7_75t_R n_7938 (.A(n_7796_o_0),
    .B(n_7812_o_0),
    .Y(n_7938_o_0));
 OAI311xp33_ASAP7_75t_R n_7939 (.A1(n_7786_o_0),
    .A2(n_7796_o_0),
    .A3(net96),
    .B1(n_7818_o_0),
    .C1(n_7938_o_0),
    .Y(n_7939_o_0));
 AOI31xp33_ASAP7_75t_R n_7940 (.A1(n_7937_o_0),
    .A2(n_7939_o_0),
    .A3(n_7916_o_0),
    .B(n_7910_o_0),
    .Y(n_7940_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7941 (.A1(n_7722_o_0),
    .A2(n_7936_o_0),
    .B(n_7940_o_0),
    .C(n_7855_o_0),
    .Y(n_7941_o_0));
 OAI21xp33_ASAP7_75t_R n_7942 (.A1(n_7822_o_0),
    .A2(n_7933_o_0),
    .B(n_7941_o_0),
    .Y(n_7942_o_0));
 OAI21xp33_ASAP7_75t_R n_7943 (.A1(n_7860_o_0),
    .A2(n_7926_o_0),
    .B(n_7942_o_0),
    .Y(n_7943_o_0));
 NAND2xp33_ASAP7_75t_R n_7944 (.A(n_7796_o_0),
    .B(n_7792_o_0),
    .Y(n_7944_o_0));
 AOI21xp33_ASAP7_75t_R n_7945 (.A1(n_7780_o_0),
    .A2(n_7796_o_0),
    .B(n_7863_o_0),
    .Y(n_7945_o_0));
 AOI211xp5_ASAP7_75t_R n_7946 (.A1(n_7944_o_0),
    .A2(n_7886_o_0),
    .B(n_7945_o_0),
    .C(n_7823_o_0),
    .Y(n_7946_o_0));
 NOR2xp33_ASAP7_75t_R n_7947 (.A(n_7796_o_0),
    .B(n_7812_o_0),
    .Y(n_7947_o_0));
 NOR3xp33_ASAP7_75t_R n_7948 (.A(n_7947_o_0),
    .B(n_7813_o_0),
    .C(n_7809_o_0),
    .Y(n_7948_o_0));
 NOR3xp33_ASAP7_75t_R n_7949 (.A(n_7948_o_0),
    .B(n_7914_o_0),
    .C(n_7714_o_0),
    .Y(n_7949_o_0));
 AOI211xp5_ASAP7_75t_R n_7950 (.A1(n_7782_o_0),
    .A2(net97),
    .B(n_7796_o_0),
    .C(n_7740_o_0),
    .Y(n_7950_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7951 (.A1(n_7740_o_0),
    .A2(n_7843_o_0),
    .B(n_7915_o_0),
    .C(n_7950_o_0),
    .Y(n_7951_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7952 (.A1(net97),
    .A2(n_7782_o_0),
    .B(n_7755_o_0),
    .C(n_7818_o_0),
    .Y(n_7952_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7953 (.A1(n_7755_o_0),
    .A2(n_7780_o_0),
    .B(n_7952_o_0),
    .C(n_7822_o_0),
    .Y(n_7953_o_0));
 AOI321xp33_ASAP7_75t_R n_7954 (.A1(n_7822_o_0),
    .A2(n_7951_o_0),
    .A3(n_7793_o_0),
    .B1(n_7935_o_0),
    .B2(n_7953_o_0),
    .C(n_7723_o_0),
    .Y(n_7954_o_0));
 INVx1_ASAP7_75t_R n_7955 (.A(n_7954_o_0),
    .Y(n_7955_o_0));
 OAI31xp33_ASAP7_75t_R n_7956 (.A1(n_7916_o_0),
    .A2(n_7946_o_0),
    .A3(n_7949_o_0),
    .B(n_7955_o_0),
    .Y(n_7956_o_0));
 NAND2xp33_ASAP7_75t_R n_7957 (.A(n_7796_o_0),
    .B(net34),
    .Y(n_7957_o_0));
 OAI31xp33_ASAP7_75t_R n_7958 (.A1(n_7782_o_0),
    .A2(n_7796_o_0),
    .A3(net97),
    .B(n_7786_o_0),
    .Y(n_7958_o_0));
 NOR2xp33_ASAP7_75t_R n_7959 (.A(n_7799_o_0),
    .B(n_7958_o_0),
    .Y(n_7959_o_0));
 AOI31xp33_ASAP7_75t_R n_7960 (.A1(n_7818_o_0),
    .A2(n_7823_o_0),
    .A3(n_7957_o_0),
    .B(n_7959_o_0),
    .Y(n_7960_o_0));
 INVx1_ASAP7_75t_R n_7961 (.A(n_7886_o_0),
    .Y(n_7961_o_0));
 INVx1_ASAP7_75t_R n_7962 (.A(n_7944_o_0),
    .Y(n_7962_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7963 (.A1(net34),
    .A2(n_7755_o_0),
    .B(n_7864_o_0),
    .C(n_7714_o_0),
    .Y(n_7963_o_0));
 OAI21xp33_ASAP7_75t_R n_7964 (.A1(n_7961_o_0),
    .A2(n_7962_o_0),
    .B(n_7963_o_0),
    .Y(n_7964_o_0));
 NAND2xp33_ASAP7_75t_R n_7965 (.A(n_7755_o_0),
    .B(n_7782_o_0),
    .Y(n_7965_o_0));
 AOI21xp33_ASAP7_75t_R n_7966 (.A1(n_7796_o_0),
    .A2(n_7780_o_0),
    .B(n_7818_o_0),
    .Y(n_7966_o_0));
 NAND2xp33_ASAP7_75t_R n_7967 (.A(n_7965_o_0),
    .B(n_7966_o_0),
    .Y(n_7967_o_0));
 AOI31xp33_ASAP7_75t_R n_7968 (.A1(n_7796_o_0),
    .A2(n_7782_o_0),
    .A3(net96),
    .B(n_7740_o_0),
    .Y(n_7968_o_0));
 OAI21xp33_ASAP7_75t_R n_7969 (.A1(n_7796_o_0),
    .A2(n_7812_o_0),
    .B(n_7968_o_0),
    .Y(n_7969_o_0));
 AOI31xp33_ASAP7_75t_R n_7970 (.A1(n_7714_o_0),
    .A2(n_7967_o_0),
    .A3(n_7969_o_0),
    .B(n_7837_o_0),
    .Y(n_7970_o_0));
 AOI21xp33_ASAP7_75t_R n_7971 (.A1(n_7964_o_0),
    .A2(n_7970_o_0),
    .B(n_7860_o_0),
    .Y(n_7971_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7972 (.A1(n_7916_o_0),
    .A2(n_7960_o_0),
    .B(n_7971_o_0),
    .C(n_7906_o_0),
    .Y(n_7972_o_0));
 OAI21xp33_ASAP7_75t_R n_7973 (.A1(n_7855_o_0),
    .A2(n_7956_o_0),
    .B(n_7972_o_0),
    .Y(n_7973_o_0));
 OAI21xp33_ASAP7_75t_R n_7974 (.A1(n_7703_o_0),
    .A2(n_7943_o_0),
    .B(n_7973_o_0),
    .Y(n_7974_o_0));
 INVx1_ASAP7_75t_R n_7975 (.A(n_7703_o_0),
    .Y(n_7975_o_0));
 INVx1_ASAP7_75t_R n_7976 (.A(n_7843_o_0),
    .Y(n_7976_o_0));
 AOI211xp5_ASAP7_75t_R n_7977 (.A1(n_7782_o_0),
    .A2(n_7755_o_0),
    .B(n_7962_o_0),
    .C(n_7786_o_0),
    .Y(n_7977_o_0));
 AOI21xp33_ASAP7_75t_R n_7978 (.A1(n_7803_o_0),
    .A2(n_7976_o_0),
    .B(n_7977_o_0),
    .Y(n_7978_o_0));
 NOR2xp33_ASAP7_75t_R n_7979 (.A(n_7879_o_0),
    .B(n_7880_o_0),
    .Y(n_7979_o_0));
 OAI31xp33_ASAP7_75t_R n_7980 (.A1(n_7818_o_0),
    .A2(n_7796_o_0),
    .A3(net34),
    .B(n_7837_o_0),
    .Y(n_7980_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_7981 (.A1(n_7783_o_0),
    .A2(n_7796_o_0),
    .B(n_7979_o_0),
    .C(n_7980_o_0),
    .Y(n_7981_o_0));
 AOI211xp5_ASAP7_75t_R n_7982 (.A1(n_7722_o_0),
    .A2(n_7978_o_0),
    .B(n_7981_o_0),
    .C(n_7823_o_0),
    .Y(n_7982_o_0));
 NOR2xp33_ASAP7_75t_R n_7983 (.A(n_7796_o_0),
    .B(n_7830_o_0),
    .Y(n_7983_o_0));
 OAI21xp33_ASAP7_75t_R n_7984 (.A1(n_7780_o_0),
    .A2(n_7755_o_0),
    .B(n_7803_o_0),
    .Y(n_7984_o_0));
 OAI31xp33_ASAP7_75t_R n_7985 (.A1(n_7740_o_0),
    .A2(n_7843_o_0),
    .A3(n_7983_o_0),
    .B(n_7984_o_0),
    .Y(n_7985_o_0));
 AOI21xp33_ASAP7_75t_R n_7986 (.A1(n_7782_o_0),
    .A2(net34),
    .B(n_7786_o_0),
    .Y(n_7986_o_0));
 OAI21xp33_ASAP7_75t_R n_7987 (.A1(net34),
    .A2(n_7796_o_0),
    .B(n_7986_o_0),
    .Y(n_7987_o_0));
 AOI21xp33_ASAP7_75t_R n_7988 (.A1(n_7786_o_0),
    .A2(n_7957_o_0),
    .B(n_7722_o_0),
    .Y(n_7988_o_0));
 AO21x1_ASAP7_75t_R n_7989 (.A1(n_7987_o_0),
    .A2(n_7988_o_0),
    .B(n_7714_o_0),
    .Y(n_7989_o_0));
 AOI21xp33_ASAP7_75t_R n_7990 (.A1(n_7722_o_0),
    .A2(n_7985_o_0),
    .B(n_7989_o_0),
    .Y(n_7990_o_0));
 AOI21xp33_ASAP7_75t_R n_7991 (.A1(n_7755_o_0),
    .A2(n_7768_o_0),
    .B(n_7740_o_0),
    .Y(n_7991_o_0));
 NAND2xp33_ASAP7_75t_R n_7992 (.A(n_7796_o_0),
    .B(n_7890_o_0),
    .Y(n_7992_o_0));
 AOI21xp33_ASAP7_75t_R n_7993 (.A1(n_7991_o_0),
    .A2(n_7992_o_0),
    .B(n_7823_o_0),
    .Y(n_7993_o_0));
 OA21x2_ASAP7_75t_R n_7994 (.A1(n_7799_o_0),
    .A2(n_7958_o_0),
    .B(n_7993_o_0),
    .Y(n_7994_o_0));
 OAI31xp33_ASAP7_75t_R n_7995 (.A1(n_7755_o_0),
    .A2(n_7768_o_0),
    .A3(net97),
    .B(n_7818_o_0),
    .Y(n_7995_o_0));
 NOR2xp33_ASAP7_75t_R n_7996 (.A(n_7796_o_0),
    .B(net97),
    .Y(n_7996_o_0));
 OAI21xp33_ASAP7_75t_R n_7997 (.A1(n_7995_o_0),
    .A2(n_7996_o_0),
    .B(n_7823_o_0),
    .Y(n_7997_o_0));
 AOI21xp33_ASAP7_75t_R n_7998 (.A1(n_7740_o_0),
    .A2(n_7920_o_0),
    .B(n_7997_o_0),
    .Y(n_7998_o_0));
 OAI21xp33_ASAP7_75t_R n_7999 (.A1(n_7921_o_0),
    .A2(n_7889_o_0),
    .B(n_7822_o_0),
    .Y(n_7999_o_0));
 INVx1_ASAP7_75t_R n_8000 (.A(n_7876_o_0),
    .Y(n_8000_o_0));
 INVx1_ASAP7_75t_R n_8001 (.A(n_7893_o_0),
    .Y(n_8001_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8002 (.A1(n_7755_o_0),
    .A2(net96),
    .B(n_7740_o_0),
    .C(n_8001_o_0),
    .Y(n_8002_o_0));
 OAI22xp33_ASAP7_75t_R n_8003 (.A1(n_7999_o_0),
    .A2(n_8000_o_0),
    .B1(n_8002_o_0),
    .B2(n_7714_o_0),
    .Y(n_8003_o_0));
 OAI321xp33_ASAP7_75t_R n_8004 (.A1(n_7837_o_0),
    .A2(n_7994_o_0),
    .A3(n_7998_o_0),
    .B1(n_8003_o_0),
    .B2(n_7722_o_0),
    .C(n_7855_o_0),
    .Y(n_8004_o_0));
 OAI31xp33_ASAP7_75t_R n_8005 (.A1(n_7708_o_0),
    .A2(n_7982_o_0),
    .A3(n_7990_o_0),
    .B(n_8004_o_0),
    .Y(n_8005_o_0));
 AOI21xp33_ASAP7_75t_R n_8006 (.A1(n_7755_o_0),
    .A2(n_7783_o_0),
    .B(n_7818_o_0),
    .Y(n_8006_o_0));
 OAI21xp33_ASAP7_75t_R n_8007 (.A1(n_7755_o_0),
    .A2(n_7890_o_0),
    .B(n_8006_o_0),
    .Y(n_8007_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8008 (.A1(n_7995_o_0),
    .A2(n_7996_o_0),
    .B(n_8007_o_0),
    .C(n_7837_o_0),
    .Y(n_8008_o_0));
 INVx1_ASAP7_75t_R n_8009 (.A(n_8008_o_0),
    .Y(n_8009_o_0));
 NOR2xp33_ASAP7_75t_R n_8010 (.A(n_7740_o_0),
    .B(n_7884_o_0),
    .Y(n_8010_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8011 (.A1(n_7796_o_0),
    .A2(n_7827_o_0),
    .B(n_8010_o_0),
    .C(n_7722_o_0),
    .Y(n_8011_o_0));
 OAI21xp33_ASAP7_75t_R n_8012 (.A1(n_7843_o_0),
    .A2(n_7802_o_0),
    .B(n_8011_o_0),
    .Y(n_8012_o_0));
 OAI211xp5_ASAP7_75t_R n_8013 (.A1(n_7832_o_0),
    .A2(n_7755_o_0),
    .B(n_7865_o_0),
    .C(n_7818_o_0),
    .Y(n_8013_o_0));
 NAND2xp33_ASAP7_75t_R n_8014 (.A(n_7796_o_0),
    .B(n_7792_o_0),
    .Y(n_8014_o_0));
 AOI31xp33_ASAP7_75t_R n_8015 (.A1(n_7786_o_0),
    .A2(n_7934_o_0),
    .A3(n_8014_o_0),
    .B(n_7837_o_0),
    .Y(n_8015_o_0));
 INVx1_ASAP7_75t_R n_8016 (.A(n_7897_o_0),
    .Y(n_8016_o_0));
 OAI211xp5_ASAP7_75t_R n_8017 (.A1(n_7812_o_0),
    .A2(n_7755_o_0),
    .B(n_7818_o_0),
    .C(n_8016_o_0),
    .Y(n_8017_o_0));
 AOI21xp33_ASAP7_75t_R n_8018 (.A1(n_8017_o_0),
    .A2(n_8001_o_0),
    .B(n_7916_o_0),
    .Y(n_8018_o_0));
 AOI211xp5_ASAP7_75t_R n_8019 (.A1(n_8013_o_0),
    .A2(n_8015_o_0),
    .B(n_8018_o_0),
    .C(n_7910_o_0),
    .Y(n_8019_o_0));
 AOI31xp33_ASAP7_75t_R n_8020 (.A1(n_7823_o_0),
    .A2(n_8009_o_0),
    .A3(n_8012_o_0),
    .B(n_8019_o_0),
    .Y(n_8020_o_0));
 NAND3xp33_ASAP7_75t_R n_8021 (.A(n_7768_o_0),
    .B(net97),
    .C(n_7755_o_0),
    .Y(n_8021_o_0));
 NAND3xp33_ASAP7_75t_R n_8022 (.A(n_8021_o_0),
    .B(n_8014_o_0),
    .C(n_7818_o_0),
    .Y(n_8022_o_0));
 AOI21xp33_ASAP7_75t_R n_8023 (.A1(n_7864_o_0),
    .A2(n_7992_o_0),
    .B(n_7837_o_0),
    .Y(n_8023_o_0));
 OAI211xp5_ASAP7_75t_R n_8024 (.A1(n_7755_o_0),
    .A2(n_7830_o_0),
    .B(n_7892_o_0),
    .C(n_7786_o_0),
    .Y(n_8024_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8025 (.A1(n_7843_o_0),
    .A2(n_7889_o_0),
    .B(n_8024_o_0),
    .C(n_7722_o_0),
    .Y(n_8025_o_0));
 AOI211xp5_ASAP7_75t_R n_8026 (.A1(n_8022_o_0),
    .A2(n_8023_o_0),
    .B(n_8025_o_0),
    .C(n_7910_o_0),
    .Y(n_8026_o_0));
 OAI211xp5_ASAP7_75t_R n_8027 (.A1(n_7812_o_0),
    .A2(n_7755_o_0),
    .B(n_7786_o_0),
    .C(n_8021_o_0),
    .Y(n_8027_o_0));
 OAI31xp33_ASAP7_75t_R n_8028 (.A1(n_7740_o_0),
    .A2(n_7866_o_0),
    .A3(n_7884_o_0),
    .B(n_8027_o_0),
    .Y(n_8028_o_0));
 AOI21xp33_ASAP7_75t_R n_8029 (.A1(n_7796_o_0),
    .A2(n_7768_o_0),
    .B(net34),
    .Y(n_8029_o_0));
 OAI22xp33_ASAP7_75t_R n_8030 (.A1(n_7783_o_0),
    .A2(n_7821_o_0),
    .B1(n_7798_o_0),
    .B2(n_7807_o_0),
    .Y(n_8030_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8031 (.A1(n_7818_o_0),
    .A2(n_8029_o_0),
    .B(n_8030_o_0),
    .C(n_7837_o_0),
    .D(n_7822_o_0),
    .Y(n_8031_o_0));
 OA21x2_ASAP7_75t_R n_8032 (.A1(n_8028_o_0),
    .A2(n_7837_o_0),
    .B(n_8031_o_0),
    .Y(n_8032_o_0));
 OAI31xp33_ASAP7_75t_R n_8033 (.A1(n_7855_o_0),
    .A2(n_8026_o_0),
    .A3(n_8032_o_0),
    .B(n_7905_o_0),
    .Y(n_8033_o_0));
 AOI21xp33_ASAP7_75t_R n_8034 (.A1(n_7708_o_0),
    .A2(n_8020_o_0),
    .B(n_8033_o_0),
    .Y(n_8034_o_0));
 AOI21xp33_ASAP7_75t_R n_8035 (.A1(n_7975_o_0),
    .A2(n_8005_o_0),
    .B(n_8034_o_0),
    .Y(n_8035_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8036 (.A1(n_7802_o_0),
    .A2(n_7861_o_0),
    .B(n_7852_o_0),
    .C(n_7722_o_0),
    .Y(n_8036_o_0));
 INVx1_ASAP7_75t_R n_8037 (.A(n_8036_o_0),
    .Y(n_8037_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8038 (.A1(n_7830_o_0),
    .A2(n_7755_o_0),
    .B(n_7813_o_0),
    .C(n_7809_o_0),
    .Y(n_8038_o_0));
 INVx1_ASAP7_75t_R n_8039 (.A(n_8038_o_0),
    .Y(n_8039_o_0));
 AOI21xp33_ASAP7_75t_R n_8040 (.A1(n_7796_o_0),
    .A2(n_7812_o_0),
    .B(n_7872_o_0),
    .Y(n_8040_o_0));
 OAI21xp33_ASAP7_75t_R n_8041 (.A1(n_8039_o_0),
    .A2(n_8040_o_0),
    .B(n_7916_o_0),
    .Y(n_8041_o_0));
 OAI21xp33_ASAP7_75t_R n_8042 (.A1(n_7755_o_0),
    .A2(n_7830_o_0),
    .B(n_7991_o_0),
    .Y(n_8042_o_0));
 OAI31xp33_ASAP7_75t_R n_8043 (.A1(n_7809_o_0),
    .A2(n_7947_o_0),
    .A3(n_7799_o_0),
    .B(n_8042_o_0),
    .Y(n_8043_o_0));
 AOI211xp5_ASAP7_75t_R n_8044 (.A1(n_8043_o_0),
    .A2(n_7837_o_0),
    .B(n_7714_o_0),
    .C(n_8023_o_0),
    .Y(n_8044_o_0));
 AOI31xp33_ASAP7_75t_R n_8045 (.A1(n_7714_o_0),
    .A2(n_8037_o_0),
    .A3(n_8041_o_0),
    .B(n_8044_o_0),
    .Y(n_8045_o_0));
 AOI21xp33_ASAP7_75t_R n_8046 (.A1(n_7850_o_0),
    .A2(n_7862_o_0),
    .B(n_7818_o_0),
    .Y(n_8046_o_0));
 INVx1_ASAP7_75t_R n_8047 (.A(n_8046_o_0),
    .Y(n_8047_o_0));
 INVx1_ASAP7_75t_R n_8048 (.A(n_7898_o_0),
    .Y(n_8048_o_0));
 NAND2xp33_ASAP7_75t_R n_8049 (.A(n_7796_o_0),
    .B(n_7798_o_0),
    .Y(n_8049_o_0));
 NAND3xp33_ASAP7_75t_R n_8050 (.A(n_8049_o_0),
    .B(n_7934_o_0),
    .C(n_7786_o_0),
    .Y(n_8050_o_0));
 OAI31xp33_ASAP7_75t_R n_8051 (.A1(n_7740_o_0),
    .A2(n_8048_o_0),
    .A3(n_7891_o_0),
    .B(n_8050_o_0),
    .Y(n_8051_o_0));
 AOI21xp33_ASAP7_75t_R n_8052 (.A1(n_7722_o_0),
    .A2(n_8051_o_0),
    .B(n_7714_o_0),
    .Y(n_8052_o_0));
 INVx1_ASAP7_75t_R n_8053 (.A(n_7872_o_0),
    .Y(n_8053_o_0));
 OAI21xp33_ASAP7_75t_R n_8054 (.A1(n_7755_o_0),
    .A2(n_7830_o_0),
    .B(n_8053_o_0),
    .Y(n_8054_o_0));
 OAI21xp33_ASAP7_75t_R n_8055 (.A1(n_7796_o_0),
    .A2(n_7798_o_0),
    .B(n_7968_o_0),
    .Y(n_8055_o_0));
 OAI21xp33_ASAP7_75t_R n_8056 (.A1(n_7958_o_0),
    .A2(n_7928_o_0),
    .B(n_8055_o_0),
    .Y(n_8056_o_0));
 AOI211xp5_ASAP7_75t_R n_8057 (.A1(_00868_),
    .A2(n_7766_o_0),
    .B(n_7792_o_0),
    .C(n_7767_o_0),
    .Y(n_8057_o_0));
 OAI21xp33_ASAP7_75t_R n_8058 (.A1(n_7842_o_0),
    .A2(n_8057_o_0),
    .B(n_7796_o_0),
    .Y(n_8058_o_0));
 AOI31xp33_ASAP7_75t_R n_8059 (.A1(n_7755_o_0),
    .A2(net96),
    .A3(n_7768_o_0),
    .B(n_7809_o_0),
    .Y(n_8059_o_0));
 AOI21xp33_ASAP7_75t_R n_8060 (.A1(n_7755_o_0),
    .A2(n_7830_o_0),
    .B(n_7995_o_0),
    .Y(n_8060_o_0));
 OAI211xp5_ASAP7_75t_R n_8061 (.A1(n_7835_o_0),
    .A2(n_7720_o_0),
    .B(n_7822_o_0),
    .C(n_7836_o_0),
    .Y(n_8061_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8062 (.A1(n_8058_o_0),
    .A2(n_8059_o_0),
    .B(n_8060_o_0),
    .C(n_8061_o_0),
    .Y(n_8062_o_0));
 OAI21xp33_ASAP7_75t_R n_8063 (.A1(n_7822_o_0),
    .A2(n_8056_o_0),
    .B(n_8062_o_0),
    .Y(n_8063_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8064 (.A1(n_8054_o_0),
    .A2(n_7867_o_0),
    .B(n_8063_o_0),
    .C(n_7975_o_0),
    .Y(n_8064_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8065 (.A1(n_8047_o_0),
    .A2(n_7995_o_0),
    .B(n_7722_o_0),
    .C(n_8052_o_0),
    .D(n_8064_o_0),
    .Y(n_8065_o_0));
 AOI21xp33_ASAP7_75t_R n_8066 (.A1(n_8045_o_0),
    .A2(n_7905_o_0),
    .B(n_8065_o_0),
    .Y(n_8066_o_0));
 OAI211xp5_ASAP7_75t_R n_8067 (.A1(n_7830_o_0),
    .A2(n_7796_o_0),
    .B(n_7786_o_0),
    .C(n_7850_o_0),
    .Y(n_8067_o_0));
 OAI31xp33_ASAP7_75t_R n_8068 (.A1(n_7740_o_0),
    .A2(n_7849_o_0),
    .A3(n_7928_o_0),
    .B(n_8067_o_0),
    .Y(n_8068_o_0));
 INVx1_ASAP7_75t_R n_8069 (.A(n_7911_o_0),
    .Y(n_8069_o_0));
 INVx1_ASAP7_75t_R n_8070 (.A(n_7801_o_0),
    .Y(n_8070_o_0));
 OAI21xp33_ASAP7_75t_R n_8071 (.A1(n_8069_o_0),
    .A2(n_8070_o_0),
    .B(n_7963_o_0),
    .Y(n_8071_o_0));
 OAI21xp33_ASAP7_75t_R n_8072 (.A1(n_7823_o_0),
    .A2(n_8068_o_0),
    .B(n_8071_o_0),
    .Y(n_8072_o_0));
 AOI211xp5_ASAP7_75t_R n_8073 (.A1(n_7801_o_0),
    .A2(n_7755_o_0),
    .B(n_7786_o_0),
    .C(n_7962_o_0),
    .Y(n_8073_o_0));
 OAI21xp33_ASAP7_75t_R n_8074 (.A1(n_8073_o_0),
    .A2(n_8046_o_0),
    .B(n_7910_o_0),
    .Y(n_8074_o_0));
 OAI311xp33_ASAP7_75t_R n_8075 (.A1(n_7796_o_0),
    .A2(n_8057_o_0),
    .A3(n_7842_o_0),
    .B1(n_7786_o_0),
    .C1(n_8014_o_0),
    .Y(n_8075_o_0));
 OAI31xp33_ASAP7_75t_R n_8076 (.A1(n_7740_o_0),
    .A2(n_7897_o_0),
    .A3(n_7921_o_0),
    .B(n_8075_o_0),
    .Y(n_8076_o_0));
 AOI21xp33_ASAP7_75t_R n_8077 (.A1(n_7714_o_0),
    .A2(n_8076_o_0),
    .B(n_7722_o_0),
    .Y(n_8077_o_0));
 AOI21xp33_ASAP7_75t_R n_8078 (.A1(n_8074_o_0),
    .A2(n_8077_o_0),
    .B(n_7905_o_0),
    .Y(n_8078_o_0));
 OAI21xp33_ASAP7_75t_R n_8079 (.A1(n_7723_o_0),
    .A2(n_8072_o_0),
    .B(n_8078_o_0),
    .Y(n_8079_o_0));
 NAND2xp33_ASAP7_75t_R n_8080 (.A(n_7991_o_0),
    .B(n_7938_o_0),
    .Y(n_8080_o_0));
 OAI31xp33_ASAP7_75t_R n_8081 (.A1(n_7842_o_0),
    .A2(n_8057_o_0),
    .A3(n_7818_o_0),
    .B(n_7755_o_0),
    .Y(n_8081_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8082 (.A1(n_7740_o_0),
    .A2(n_7768_o_0),
    .B(n_7755_o_0),
    .C(n_8081_o_0),
    .Y(n_8082_o_0));
 OAI21xp33_ASAP7_75t_R n_8083 (.A1(n_7786_o_0),
    .A2(n_8021_o_0),
    .B(n_7714_o_0),
    .Y(n_8083_o_0));
 AOI31xp33_ASAP7_75t_R n_8084 (.A1(n_7786_o_0),
    .A2(n_7892_o_0),
    .A3(n_8049_o_0),
    .B(n_8083_o_0),
    .Y(n_8084_o_0));
 AOI31xp33_ASAP7_75t_R n_8085 (.A1(n_7823_o_0),
    .A2(n_8080_o_0),
    .A3(n_8082_o_0),
    .B(n_8084_o_0),
    .Y(n_8085_o_0));
 INVx1_ASAP7_75t_R n_8086 (.A(n_7833_o_0),
    .Y(n_8086_o_0));
 OAI21xp33_ASAP7_75t_R n_8087 (.A1(n_7842_o_0),
    .A2(n_8057_o_0),
    .B(n_7911_o_0),
    .Y(n_8087_o_0));
 OAI31xp33_ASAP7_75t_R n_8088 (.A1(n_7809_o_0),
    .A2(n_7799_o_0),
    .A3(n_7996_o_0),
    .B(n_8087_o_0),
    .Y(n_8088_o_0));
 AND4x1_ASAP7_75t_R n_8089 (.A(n_7801_o_0),
    .B(n_7786_o_0),
    .C(n_7755_o_0),
    .D(n_7714_o_0),
    .Y(n_8089_o_0));
 AOI21xp33_ASAP7_75t_R n_8090 (.A1(n_7823_o_0),
    .A2(n_8088_o_0),
    .B(n_8089_o_0),
    .Y(n_8090_o_0));
 AOI21xp33_ASAP7_75t_R n_8091 (.A1(n_8086_o_0),
    .A2(n_8090_o_0),
    .B(n_7975_o_0),
    .Y(n_8091_o_0));
 OAI21xp33_ASAP7_75t_R n_8092 (.A1(n_7916_o_0),
    .A2(n_8085_o_0),
    .B(n_8091_o_0),
    .Y(n_8092_o_0));
 AO21x1_ASAP7_75t_R n_8093 (.A1(n_8079_o_0),
    .A2(n_8092_o_0),
    .B(n_7860_o_0),
    .Y(n_8093_o_0));
 OAI21xp33_ASAP7_75t_R n_8094 (.A1(n_7708_o_0),
    .A2(n_8066_o_0),
    .B(n_8093_o_0),
    .Y(n_8094_o_0));
 OAI21xp33_ASAP7_75t_R n_8095 (.A1(n_7755_o_0),
    .A2(n_7782_o_0),
    .B(net34),
    .Y(n_8095_o_0));
 AOI21xp33_ASAP7_75t_R n_8096 (.A1(n_7898_o_0),
    .A2(n_7927_o_0),
    .B(n_7818_o_0),
    .Y(n_8096_o_0));
 INVx1_ASAP7_75t_R n_8097 (.A(n_8096_o_0),
    .Y(n_8097_o_0));
 OAI211xp5_ASAP7_75t_R n_8098 (.A1(n_8095_o_0),
    .A2(n_7740_o_0),
    .B(n_8097_o_0),
    .C(n_7916_o_0),
    .Y(n_8098_o_0));
 OAI21xp33_ASAP7_75t_R n_8099 (.A1(net34),
    .A2(n_7755_o_0),
    .B(n_7864_o_0),
    .Y(n_8099_o_0));
 OAI31xp33_ASAP7_75t_R n_8100 (.A1(n_7740_o_0),
    .A2(n_7861_o_0),
    .A3(n_7996_o_0),
    .B(n_8099_o_0),
    .Y(n_8100_o_0));
 AOI21xp33_ASAP7_75t_R n_8101 (.A1(n_7837_o_0),
    .A2(n_8100_o_0),
    .B(n_7855_o_0),
    .Y(n_8101_o_0));
 OAI211xp5_ASAP7_75t_R n_8102 (.A1(n_7783_o_0),
    .A2(n_7796_o_0),
    .B(n_7944_o_0),
    .C(n_7809_o_0),
    .Y(n_8102_o_0));
 NOR2xp33_ASAP7_75t_R n_8103 (.A(n_7755_o_0),
    .B(net97),
    .Y(n_8103_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8104 (.A1(n_7849_o_0),
    .A2(n_8103_o_0),
    .B(n_7809_o_0),
    .C(n_7847_o_0),
    .Y(n_8104_o_0));
 AOI31xp33_ASAP7_75t_R n_8105 (.A1(n_7722_o_0),
    .A2(n_8007_o_0),
    .A3(n_8102_o_0),
    .B(n_8104_o_0),
    .Y(n_8105_o_0));
 OAI21xp33_ASAP7_75t_R n_8106 (.A1(n_7856_o_0),
    .A2(n_8105_o_0),
    .B(n_7910_o_0),
    .Y(n_8106_o_0));
 INVx1_ASAP7_75t_R n_8107 (.A(n_7952_o_0),
    .Y(n_8107_o_0));
 AOI21xp33_ASAP7_75t_R n_8108 (.A1(n_7796_o_0),
    .A2(n_7801_o_0),
    .B(n_8107_o_0),
    .Y(n_8108_o_0));
 NAND2xp33_ASAP7_75t_R n_8109 (.A(n_7796_o_0),
    .B(n_7809_o_0),
    .Y(n_8109_o_0));
 OAI221xp5_ASAP7_75t_R n_8110 (.A1(n_7783_o_0),
    .A2(n_7821_o_0),
    .B1(n_7801_o_0),
    .B2(n_8109_o_0),
    .C(n_8021_o_0),
    .Y(n_8110_o_0));
 OA22x2_ASAP7_75t_R n_8111 (.A1(n_8108_o_0),
    .A2(n_7838_o_0),
    .B1(n_8110_o_0),
    .B2(n_7723_o_0),
    .Y(n_8111_o_0));
 OAI21xp33_ASAP7_75t_R n_8112 (.A1(n_7796_o_0),
    .A2(n_7832_o_0),
    .B(n_7834_o_0),
    .Y(n_8112_o_0));
 AOI21xp33_ASAP7_75t_R n_8113 (.A1(n_7916_o_0),
    .A2(n_8112_o_0),
    .B(n_7708_o_0),
    .Y(n_8113_o_0));
 NOR3xp33_ASAP7_75t_R n_8114 (.A(n_7797_o_0),
    .B(n_8103_o_0),
    .C(n_7740_o_0),
    .Y(n_8114_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8115 (.A1(n_7966_o_0),
    .A2(n_7965_o_0),
    .B(n_8114_o_0),
    .C(n_7723_o_0),
    .Y(n_8115_o_0));
 AOI21xp33_ASAP7_75t_R n_8116 (.A1(n_8113_o_0),
    .A2(n_8115_o_0),
    .B(n_7823_o_0),
    .Y(n_8116_o_0));
 OAI21xp33_ASAP7_75t_R n_8117 (.A1(n_7856_o_0),
    .A2(n_8111_o_0),
    .B(n_8116_o_0),
    .Y(n_8117_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8118 (.A1(n_8098_o_0),
    .A2(n_8101_o_0),
    .B(n_8106_o_0),
    .C(n_8117_o_0),
    .Y(n_8118_o_0));
 NAND2xp33_ASAP7_75t_R n_8119 (.A(n_7944_o_0),
    .B(n_7886_o_0),
    .Y(n_8119_o_0));
 AOI31xp33_ASAP7_75t_R n_8120 (.A1(net34),
    .A2(n_7796_o_0),
    .A3(n_7740_o_0),
    .B(n_7723_o_0),
    .Y(n_8120_o_0));
 AOI211xp5_ASAP7_75t_R n_8121 (.A1(n_7864_o_0),
    .A2(n_7938_o_0),
    .B(n_7911_o_0),
    .C(n_7916_o_0),
    .Y(n_8121_o_0));
 AOI31xp33_ASAP7_75t_R n_8122 (.A1(n_7876_o_0),
    .A2(n_8119_o_0),
    .A3(n_8120_o_0),
    .B(n_8121_o_0),
    .Y(n_8122_o_0));
 OAI21xp33_ASAP7_75t_R n_8123 (.A1(n_7861_o_0),
    .A2(n_7866_o_0),
    .B(n_7809_o_0),
    .Y(n_8123_o_0));
 INVx1_ASAP7_75t_R n_8124 (.A(n_7793_o_0),
    .Y(n_8124_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8125 (.A1(n_8124_o_0),
    .A2(n_7781_o_0),
    .B(n_7740_o_0),
    .C(n_7916_o_0),
    .Y(n_8125_o_0));
 AOI21xp33_ASAP7_75t_R n_8126 (.A1(n_8123_o_0),
    .A2(n_8125_o_0),
    .B(n_7860_o_0),
    .Y(n_8126_o_0));
 OAI211xp5_ASAP7_75t_R n_8127 (.A1(n_7866_o_0),
    .A2(n_7834_o_0),
    .B(n_8097_o_0),
    .C(n_7722_o_0),
    .Y(n_8127_o_0));
 AOI22xp33_ASAP7_75t_R n_8128 (.A1(n_8122_o_0),
    .A2(n_7856_o_0),
    .B1(n_8126_o_0),
    .B2(n_8127_o_0),
    .Y(n_8128_o_0));
 OAI21xp33_ASAP7_75t_R n_8129 (.A1(n_7796_o_0),
    .A2(n_7827_o_0),
    .B(n_7976_o_0),
    .Y(n_8129_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8130 (.A1(n_7809_o_0),
    .A2(n_8129_o_0),
    .B(n_7819_o_0),
    .C(n_7916_o_0),
    .Y(n_8130_o_0));
 OAI21xp33_ASAP7_75t_R n_8131 (.A1(n_7755_o_0),
    .A2(n_7780_o_0),
    .B(n_7740_o_0),
    .Y(n_8131_o_0));
 OAI21xp33_ASAP7_75t_R n_8132 (.A1(n_7786_o_0),
    .A2(n_7871_o_0),
    .B(n_8131_o_0),
    .Y(n_8132_o_0));
 AO21x1_ASAP7_75t_R n_8133 (.A1(n_8132_o_0),
    .A2(n_7916_o_0),
    .B(n_7708_o_0),
    .Y(n_8133_o_0));
 AOI21xp33_ASAP7_75t_R n_8134 (.A1(net34),
    .A2(n_7755_o_0),
    .B(n_7834_o_0),
    .Y(n_8134_o_0));
 OAI221xp5_ASAP7_75t_R n_8135 (.A1(n_7809_o_0),
    .A2(n_7890_o_0),
    .B1(n_7740_o_0),
    .B2(n_7843_o_0),
    .C(n_7723_o_0),
    .Y(n_8135_o_0));
 OAI31xp33_ASAP7_75t_R n_8136 (.A1(n_7723_o_0),
    .A2(n_7828_o_0),
    .A3(n_8134_o_0),
    .B(n_8135_o_0),
    .Y(n_8136_o_0));
 AOI21xp33_ASAP7_75t_R n_8137 (.A1(n_7855_o_0),
    .A2(n_8136_o_0),
    .B(n_7823_o_0),
    .Y(n_8137_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8138 (.A1(n_8130_o_0),
    .A2(n_8133_o_0),
    .B(n_8137_o_0),
    .C(n_7906_o_0),
    .Y(n_8138_o_0));
 OAI21xp33_ASAP7_75t_R n_8139 (.A1(n_7714_o_0),
    .A2(n_8128_o_0),
    .B(n_8138_o_0),
    .Y(n_8139_o_0));
 OA21x2_ASAP7_75t_R n_8140 (.A1(n_8118_o_0),
    .A2(n_7703_o_0),
    .B(n_8139_o_0),
    .Y(n_8140_o_0));
 OAI21xp33_ASAP7_75t_R n_8141 (.A1(n_7740_o_0),
    .A2(net96),
    .B(n_7822_o_0),
    .Y(n_8141_o_0));
 NAND2xp33_ASAP7_75t_R n_8142 (.A(n_7786_o_0),
    .B(n_7992_o_0),
    .Y(n_8142_o_0));
 OA21x2_ASAP7_75t_R n_8143 (.A1(n_7889_o_0),
    .A2(n_7781_o_0),
    .B(n_7910_o_0),
    .Y(n_8143_o_0));
 AOI21xp33_ASAP7_75t_R n_8144 (.A1(n_8142_o_0),
    .A2(n_8143_o_0),
    .B(n_7856_o_0),
    .Y(n_8144_o_0));
 OAI21xp33_ASAP7_75t_R n_8145 (.A1(n_7796_o_0),
    .A2(n_7827_o_0),
    .B(n_7938_o_0),
    .Y(n_8145_o_0));
 OAI21xp33_ASAP7_75t_R n_8146 (.A1(n_7740_o_0),
    .A2(n_8145_o_0),
    .B(n_7901_o_0),
    .Y(n_8146_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8147 (.A1(n_8038_o_0),
    .A2(n_7872_o_0),
    .B(n_7714_o_0),
    .C(n_7860_o_0),
    .Y(n_8147_o_0));
 AOI21xp33_ASAP7_75t_R n_8148 (.A1(n_7822_o_0),
    .A2(n_8146_o_0),
    .B(n_8147_o_0),
    .Y(n_8148_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8149 (.A1(n_8096_o_0),
    .A2(n_8141_o_0),
    .B(n_8144_o_0),
    .C(n_8148_o_0),
    .Y(n_8149_o_0));
 OAI211xp5_ASAP7_75t_R n_8150 (.A1(n_7783_o_0),
    .A2(n_7796_o_0),
    .B(n_8049_o_0),
    .C(n_7786_o_0),
    .Y(n_8150_o_0));
 OAI31xp33_ASAP7_75t_R n_8151 (.A1(n_7740_o_0),
    .A2(n_7768_o_0),
    .A3(n_7921_o_0),
    .B(n_8150_o_0),
    .Y(n_8151_o_0));
 NAND2xp33_ASAP7_75t_R n_8152 (.A(n_7714_o_0),
    .B(n_8151_o_0),
    .Y(n_8152_o_0));
 OAI21xp33_ASAP7_75t_R n_8153 (.A1(n_7921_o_0),
    .A2(n_8006_o_0),
    .B(n_7910_o_0),
    .Y(n_8153_o_0));
 NAND3xp33_ASAP7_75t_R n_8154 (.A(n_7814_o_0),
    .B(n_7927_o_0),
    .C(n_7786_o_0),
    .Y(n_8154_o_0));
 AOI21xp33_ASAP7_75t_R n_8155 (.A1(n_7755_o_0),
    .A2(n_7812_o_0),
    .B(n_7786_o_0),
    .Y(n_8155_o_0));
 OAI21xp33_ASAP7_75t_R n_8156 (.A1(n_7755_o_0),
    .A2(n_7830_o_0),
    .B(n_8155_o_0),
    .Y(n_8156_o_0));
 OAI22xp33_ASAP7_75t_R n_8157 (.A1(n_8131_o_0),
    .A2(n_7996_o_0),
    .B1(n_7801_o_0),
    .B2(n_8109_o_0),
    .Y(n_8157_o_0));
 AOI321xp33_ASAP7_75t_R n_8158 (.A1(n_8154_o_0),
    .A2(n_8156_o_0),
    .A3(n_7822_o_0),
    .B1(n_8157_o_0),
    .B2(n_7910_o_0),
    .C(n_7856_o_0),
    .Y(n_8158_o_0));
 AOI31xp33_ASAP7_75t_R n_8159 (.A1(n_7860_o_0),
    .A2(n_8152_o_0),
    .A3(n_8153_o_0),
    .B(n_8158_o_0),
    .Y(n_8159_o_0));
 AOI22xp33_ASAP7_75t_R n_8160 (.A1(n_8149_o_0),
    .A2(n_7723_o_0),
    .B1(n_7916_o_0),
    .B2(n_8159_o_0),
    .Y(n_8160_o_0));
 NOR2xp33_ASAP7_75t_R n_8161 (.A(n_7884_o_0),
    .B(n_7889_o_0),
    .Y(n_8161_o_0));
 AOI31xp33_ASAP7_75t_R n_8162 (.A1(n_7786_o_0),
    .A2(n_7898_o_0),
    .A3(n_8049_o_0),
    .B(n_8161_o_0),
    .Y(n_8162_o_0));
 OAI21xp33_ASAP7_75t_R n_8163 (.A1(n_7861_o_0),
    .A2(n_7863_o_0),
    .B(n_7723_o_0),
    .Y(n_8163_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8164 (.A1(n_7818_o_0),
    .A2(n_7768_o_0),
    .B(n_8163_o_0),
    .C(n_7714_o_0),
    .Y(n_8164_o_0));
 OAI31xp33_ASAP7_75t_R n_8165 (.A1(n_7809_o_0),
    .A2(n_7797_o_0),
    .A3(n_7921_o_0),
    .B(n_7819_o_0),
    .Y(n_8165_o_0));
 AOI21xp33_ASAP7_75t_R n_8166 (.A1(n_8059_o_0),
    .A2(n_7938_o_0),
    .B(n_7837_o_0),
    .Y(n_8166_o_0));
 OAI21xp33_ASAP7_75t_R n_8167 (.A1(n_8069_o_0),
    .A2(n_7830_o_0),
    .B(n_8166_o_0),
    .Y(n_8167_o_0));
 OAI211xp5_ASAP7_75t_R n_8168 (.A1(n_7722_o_0),
    .A2(n_8165_o_0),
    .B(n_8167_o_0),
    .C(n_7823_o_0),
    .Y(n_8168_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8169 (.A1(n_8162_o_0),
    .A2(n_7916_o_0),
    .B(n_8164_o_0),
    .C(n_8168_o_0),
    .Y(n_8169_o_0));
 AOI21xp33_ASAP7_75t_R n_8170 (.A1(n_7818_o_0),
    .A2(n_7798_o_0),
    .B(n_7722_o_0),
    .Y(n_8170_o_0));
 NAND2xp33_ASAP7_75t_R n_8171 (.A(n_7796_o_0),
    .B(n_7830_o_0),
    .Y(n_8171_o_0));
 NOR3xp33_ASAP7_75t_R n_8172 (.A(n_8057_o_0),
    .B(n_7842_o_0),
    .C(n_7796_o_0),
    .Y(n_8172_o_0));
 OAI31xp33_ASAP7_75t_R n_8173 (.A1(n_7809_o_0),
    .A2(n_7891_o_0),
    .A3(n_8172_o_0),
    .B(n_7916_o_0),
    .Y(n_8173_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8174 (.A1(n_8171_o_0),
    .A2(n_7914_o_0),
    .B(n_8173_o_0),
    .C(n_7823_o_0),
    .Y(n_8174_o_0));
 NOR2xp33_ASAP7_75t_R n_8175 (.A(n_7991_o_0),
    .B(n_7722_o_0),
    .Y(n_8175_o_0));
 OAI21xp33_ASAP7_75t_R n_8176 (.A1(n_7947_o_0),
    .A2(n_8001_o_0),
    .B(n_8175_o_0),
    .Y(n_8176_o_0));
 OAI21xp33_ASAP7_75t_R n_8177 (.A1(n_7755_o_0),
    .A2(n_7890_o_0),
    .B(n_7809_o_0),
    .Y(n_8177_o_0));
 OAI211xp5_ASAP7_75t_R n_8178 (.A1(n_7783_o_0),
    .A2(n_7821_o_0),
    .B(n_8177_o_0),
    .C(n_7722_o_0),
    .Y(n_8178_o_0));
 NAND3xp33_ASAP7_75t_R n_8179 (.A(n_8176_o_0),
    .B(n_8178_o_0),
    .C(n_7822_o_0),
    .Y(n_8179_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8180 (.A1(n_7958_o_0),
    .A2(n_8170_o_0),
    .B(n_8174_o_0),
    .C(n_8179_o_0),
    .Y(n_8180_o_0));
 OAI22xp33_ASAP7_75t_R n_8181 (.A1(n_8169_o_0),
    .A2(n_7855_o_0),
    .B1(n_7860_o_0),
    .B2(n_8180_o_0),
    .Y(n_8181_o_0));
 OAI22xp33_ASAP7_75t_R n_8182 (.A1(n_8160_o_0),
    .A2(n_7703_o_0),
    .B1(n_8181_o_0),
    .B2(n_7906_o_0),
    .Y(n_8182_o_0));
 AOI211xp5_ASAP7_75t_R n_8183 (.A1(n_7832_o_0),
    .A2(n_7796_o_0),
    .B(n_8172_o_0),
    .C(n_7809_o_0),
    .Y(n_8183_o_0));
 AOI31xp33_ASAP7_75t_R n_8184 (.A1(n_7818_o_0),
    .A2(n_7898_o_0),
    .A3(n_7885_o_0),
    .B(n_8183_o_0),
    .Y(n_8184_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8185 (.A1(n_7916_o_0),
    .A2(n_8184_o_0),
    .B(n_7822_o_0),
    .C(n_7881_o_0),
    .Y(n_8185_o_0));
 NAND2xp33_ASAP7_75t_R n_8186 (.A(n_7755_o_0),
    .B(n_7801_o_0),
    .Y(n_8186_o_0));
 OAI221xp5_ASAP7_75t_R n_8187 (.A1(n_8186_o_0),
    .A2(n_7809_o_0),
    .B1(n_7823_o_0),
    .B2(n_8002_o_0),
    .C(n_7916_o_0),
    .Y(n_8187_o_0));
 INVx1_ASAP7_75t_R n_8188 (.A(n_8187_o_0),
    .Y(n_8188_o_0));
 AOI21xp33_ASAP7_75t_R n_8189 (.A1(n_7755_o_0),
    .A2(n_7827_o_0),
    .B(n_7786_o_0),
    .Y(n_8189_o_0));
 AOI211xp5_ASAP7_75t_R n_8190 (.A1(n_7755_o_0),
    .A2(n_7768_o_0),
    .B(n_7843_o_0),
    .C(n_7809_o_0),
    .Y(n_8190_o_0));
 AOI21xp33_ASAP7_75t_R n_8191 (.A1(n_8189_o_0),
    .A2(n_7850_o_0),
    .B(n_8190_o_0),
    .Y(n_8191_o_0));
 OAI21xp33_ASAP7_75t_R n_8192 (.A1(net34),
    .A2(n_7755_o_0),
    .B(n_8189_o_0),
    .Y(n_8192_o_0));
 OAI31xp33_ASAP7_75t_R n_8193 (.A1(n_7809_o_0),
    .A2(n_7830_o_0),
    .A3(n_7755_o_0),
    .B(n_8192_o_0),
    .Y(n_8193_o_0));
 AOI21xp33_ASAP7_75t_R n_8194 (.A1(n_7722_o_0),
    .A2(n_8193_o_0),
    .B(n_7714_o_0),
    .Y(n_8194_o_0));
 OAI21xp33_ASAP7_75t_R n_8195 (.A1(n_7916_o_0),
    .A2(n_8191_o_0),
    .B(n_8194_o_0),
    .Y(n_8195_o_0));
 OAI211xp5_ASAP7_75t_R n_8196 (.A1(n_8185_o_0),
    .A2(n_8188_o_0),
    .B(n_7855_o_0),
    .C(n_8195_o_0),
    .Y(n_8196_o_0));
 OAI21xp33_ASAP7_75t_R n_8197 (.A1(n_7786_o_0),
    .A2(n_8021_o_0),
    .B(n_7722_o_0),
    .Y(n_8197_o_0));
 NOR2xp33_ASAP7_75t_R n_8198 (.A(n_7863_o_0),
    .B(n_7843_o_0),
    .Y(n_8198_o_0));
 NOR2xp33_ASAP7_75t_R n_8199 (.A(n_7768_o_0),
    .B(n_8069_o_0),
    .Y(n_8199_o_0));
 OAI21xp33_ASAP7_75t_R n_8200 (.A1(n_7755_o_0),
    .A2(n_7830_o_0),
    .B(n_7952_o_0),
    .Y(n_8200_o_0));
 AOI31xp33_ASAP7_75t_R n_8201 (.A1(n_7755_o_0),
    .A2(n_7809_o_0),
    .A3(n_7780_o_0),
    .B(n_7916_o_0),
    .Y(n_8201_o_0));
 OAI311xp33_ASAP7_75t_R n_8202 (.A1(n_7740_o_0),
    .A2(n_7890_o_0),
    .A3(n_7755_o_0),
    .B1(n_8200_o_0),
    .C1(n_8201_o_0),
    .Y(n_8202_o_0));
 OAI31xp33_ASAP7_75t_R n_8203 (.A1(n_8197_o_0),
    .A2(n_8198_o_0),
    .A3(n_8199_o_0),
    .B(n_8202_o_0),
    .Y(n_8203_o_0));
 NOR2xp33_ASAP7_75t_R n_8204 (.A(n_7832_o_0),
    .B(n_8109_o_0),
    .Y(n_8204_o_0));
 AO21x1_ASAP7_75t_R n_8205 (.A1(n_7927_o_0),
    .A2(n_7898_o_0),
    .B(n_7786_o_0),
    .Y(n_8205_o_0));
 OAI21xp33_ASAP7_75t_R n_8206 (.A1(net96),
    .A2(n_7818_o_0),
    .B(n_8205_o_0),
    .Y(n_8206_o_0));
 OAI32xp33_ASAP7_75t_R n_8207 (.A1(n_8000_o_0),
    .A2(n_8197_o_0),
    .A3(n_8204_o_0),
    .B1(n_8206_o_0),
    .B2(n_7916_o_0),
    .Y(n_8207_o_0));
 OAI22xp33_ASAP7_75t_R n_8208 (.A1(n_8203_o_0),
    .A2(n_7714_o_0),
    .B1(n_7823_o_0),
    .B2(n_8207_o_0),
    .Y(n_8208_o_0));
 AOI21xp33_ASAP7_75t_R n_8209 (.A1(n_7860_o_0),
    .A2(n_8208_o_0),
    .B(n_7905_o_0),
    .Y(n_8209_o_0));
 AOI21xp33_ASAP7_75t_R n_8210 (.A1(n_7796_o_0),
    .A2(n_7830_o_0),
    .B(n_7818_o_0),
    .Y(n_8210_o_0));
 OA21x2_ASAP7_75t_R n_8211 (.A1(n_8134_o_0),
    .A2(n_8210_o_0),
    .B(n_7916_o_0),
    .Y(n_8211_o_0));
 NOR2xp33_ASAP7_75t_R n_8212 (.A(n_7809_o_0),
    .B(n_8048_o_0),
    .Y(n_8212_o_0));
 XNOR2xp5_ASAP7_75t_R n_8213 (.A(n_7755_o_0),
    .B(net34),
    .Y(n_8213_o_0));
 AOI22xp33_ASAP7_75t_R n_8214 (.A1(n_8212_o_0),
    .A2(n_8049_o_0),
    .B1(n_7818_o_0),
    .B2(n_8213_o_0),
    .Y(n_8214_o_0));
 AOI22xp33_ASAP7_75t_R n_8215 (.A1(n_7914_o_0),
    .A2(n_7992_o_0),
    .B1(n_7786_o_0),
    .B2(n_7850_o_0),
    .Y(n_8215_o_0));
 AOI21xp33_ASAP7_75t_R n_8216 (.A1(n_7722_o_0),
    .A2(n_8215_o_0),
    .B(n_7823_o_0),
    .Y(n_8216_o_0));
 OAI21xp33_ASAP7_75t_R n_8217 (.A1(n_7916_o_0),
    .A2(n_8214_o_0),
    .B(n_8216_o_0),
    .Y(n_8217_o_0));
 OAI311xp33_ASAP7_75t_R n_8218 (.A1(n_7714_o_0),
    .A2(n_8211_o_0),
    .A3(n_8011_o_0),
    .B1(n_7855_o_0),
    .C1(n_8217_o_0),
    .Y(n_8218_o_0));
 NOR3xp33_ASAP7_75t_R n_8219 (.A(n_7851_o_0),
    .B(n_7861_o_0),
    .C(n_7740_o_0),
    .Y(n_8219_o_0));
 XOR2xp5_ASAP7_75t_R n_822 (.A(_00442_),
    .B(_00880_),
    .Y(n_822_o_0));
 AOI31xp33_ASAP7_75t_R n_8220 (.A1(n_7922_o_0),
    .A2(n_8212_o_0),
    .A3(n_7740_o_0),
    .B(n_8219_o_0),
    .Y(n_8220_o_0));
 OAI211xp5_ASAP7_75t_R n_8221 (.A1(n_7818_o_0),
    .A2(n_7934_o_0),
    .B(n_8038_o_0),
    .C(n_7823_o_0),
    .Y(n_8221_o_0));
 OAI21xp33_ASAP7_75t_R n_8222 (.A1(n_7910_o_0),
    .A2(n_8220_o_0),
    .B(n_8221_o_0),
    .Y(n_8222_o_0));
 OAI22xp33_ASAP7_75t_R n_8223 (.A1(n_8001_o_0),
    .A2(n_7797_o_0),
    .B1(n_7740_o_0),
    .B2(n_7920_o_0),
    .Y(n_8223_o_0));
 OAI21xp33_ASAP7_75t_R n_8224 (.A1(n_7952_o_0),
    .A2(n_7986_o_0),
    .B(n_7822_o_0),
    .Y(n_8224_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8225 (.A1(n_7768_o_0),
    .A2(n_7796_o_0),
    .B(n_8224_o_0),
    .C(n_7722_o_0),
    .Y(n_8225_o_0));
 AOI21xp33_ASAP7_75t_R n_8226 (.A1(n_7910_o_0),
    .A2(n_8223_o_0),
    .B(n_8225_o_0),
    .Y(n_8226_o_0));
 AOI21xp33_ASAP7_75t_R n_8227 (.A1(n_7837_o_0),
    .A2(n_8222_o_0),
    .B(n_8226_o_0),
    .Y(n_8227_o_0));
 AOI21xp33_ASAP7_75t_R n_8228 (.A1(n_7860_o_0),
    .A2(n_8227_o_0),
    .B(n_7975_o_0),
    .Y(n_8228_o_0));
 AOI22xp33_ASAP7_75t_R n_8229 (.A1(n_8196_o_0),
    .A2(n_8209_o_0),
    .B1(n_8218_o_0),
    .B2(n_8228_o_0),
    .Y(n_8229_o_0));
 XNOR2xp5_ASAP7_75t_R n_823 (.A(_00912_),
    .B(n_822_o_0),
    .Y(n_823_o_0));
 AOI31xp33_ASAP7_75t_R n_8230 (.A1(n_7786_o_0),
    .A2(n_7992_o_0),
    .A3(n_7934_o_0),
    .B(n_8189_o_0),
    .Y(n_8230_o_0));
 OAI21xp33_ASAP7_75t_R n_8231 (.A1(n_7723_o_0),
    .A2(n_8230_o_0),
    .B(n_7910_o_0),
    .Y(n_8231_o_0));
 NOR3xp33_ASAP7_75t_R n_8232 (.A(n_8053_o_0),
    .B(n_8155_o_0),
    .C(n_7916_o_0),
    .Y(n_8232_o_0));
 OAI21xp33_ASAP7_75t_R n_8233 (.A1(n_7768_o_0),
    .A2(n_7818_o_0),
    .B(n_7722_o_0),
    .Y(n_8233_o_0));
 OAI311xp33_ASAP7_75t_R n_8234 (.A1(n_7782_o_0),
    .A2(net34),
    .A3(n_7755_o_0),
    .B1(n_7786_o_0),
    .C1(n_7898_o_0),
    .Y(n_8234_o_0));
 OAI31xp33_ASAP7_75t_R n_8235 (.A1(n_7740_o_0),
    .A2(n_7861_o_0),
    .A3(n_7996_o_0),
    .B(n_8234_o_0),
    .Y(n_8235_o_0));
 AOI21xp33_ASAP7_75t_R n_8236 (.A1(n_7837_o_0),
    .A2(n_8235_o_0),
    .B(n_7823_o_0),
    .Y(n_8236_o_0));
 OAI21xp33_ASAP7_75t_R n_8237 (.A1(n_8114_o_0),
    .A2(n_8233_o_0),
    .B(n_8236_o_0),
    .Y(n_8237_o_0));
 OA21x2_ASAP7_75t_R n_8238 (.A1(n_8231_o_0),
    .A2(n_8232_o_0),
    .B(n_8237_o_0),
    .Y(n_8238_o_0));
 INVx1_ASAP7_75t_R n_8239 (.A(n_8082_o_0),
    .Y(n_8239_o_0));
 XNOR2xp5_ASAP7_75t_R n_824 (.A(_00944_),
    .B(n_823_o_0),
    .Y(n_824_o_0));
 OAI21xp33_ASAP7_75t_R n_8240 (.A1(n_7919_o_0),
    .A2(n_8239_o_0),
    .B(n_7916_o_0),
    .Y(n_8240_o_0));
 INVx1_ASAP7_75t_R n_8241 (.A(n_8200_o_0),
    .Y(n_8241_o_0));
 OAI21xp33_ASAP7_75t_R n_8242 (.A1(n_7977_o_0),
    .A2(n_8241_o_0),
    .B(n_7723_o_0),
    .Y(n_8242_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8243 (.A1(net96),
    .A2(n_7796_o_0),
    .B(n_7782_o_0),
    .C(n_7809_o_0),
    .Y(n_8243_o_0));
 AOI211xp5_ASAP7_75t_R n_8244 (.A1(n_7812_o_0),
    .A2(n_7911_o_0),
    .B(n_8243_o_0),
    .C(n_7950_o_0),
    .Y(n_8244_o_0));
 AOI21xp33_ASAP7_75t_R n_8245 (.A1(n_7916_o_0),
    .A2(n_8244_o_0),
    .B(n_7910_o_0),
    .Y(n_8245_o_0));
 OAI31xp33_ASAP7_75t_R n_8246 (.A1(n_7722_o_0),
    .A2(n_7952_o_0),
    .A3(n_8134_o_0),
    .B(n_8245_o_0),
    .Y(n_8246_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8247 (.A1(n_8240_o_0),
    .A2(n_8242_o_0),
    .B(n_7714_o_0),
    .C(n_8246_o_0),
    .Y(n_8247_o_0));
 OAI22xp33_ASAP7_75t_R n_8248 (.A1(n_8238_o_0),
    .A2(n_7860_o_0),
    .B1(n_7855_o_0),
    .B2(n_8247_o_0),
    .Y(n_8248_o_0));
 INVx1_ASAP7_75t_R n_8249 (.A(n_7828_o_0),
    .Y(n_8249_o_0));
 INVx1_ASAP7_75t_R n_825 (.A(_00976_),
    .Y(n_825_o_0));
 AOI321xp33_ASAP7_75t_R n_8250 (.A1(n_7780_o_0),
    .A2(n_8069_o_0),
    .A3(n_7796_o_0),
    .B1(n_7818_o_0),
    .B2(n_7812_o_0),
    .C(n_7916_o_0),
    .Y(n_8250_o_0));
 AOI31xp33_ASAP7_75t_R n_8251 (.A1(n_8249_o_0),
    .A2(n_8119_o_0),
    .A3(n_8120_o_0),
    .B(n_8250_o_0),
    .Y(n_8251_o_0));
 INVx1_ASAP7_75t_R n_8252 (.A(n_8251_o_0),
    .Y(n_8252_o_0));
 NAND3xp33_ASAP7_75t_R n_8253 (.A(n_8058_o_0),
    .B(n_8021_o_0),
    .C(n_7786_o_0),
    .Y(n_8253_o_0));
 AOI21xp33_ASAP7_75t_R n_8254 (.A1(n_7818_o_0),
    .A2(n_7957_o_0),
    .B(n_7722_o_0),
    .Y(n_8254_o_0));
 OAI21xp33_ASAP7_75t_R n_8255 (.A1(n_7996_o_0),
    .A2(n_7915_o_0),
    .B(n_7916_o_0),
    .Y(n_8255_o_0));
 AOI21xp33_ASAP7_75t_R n_8256 (.A1(n_7976_o_0),
    .A2(n_7914_o_0),
    .B(n_8255_o_0),
    .Y(n_8256_o_0));
 AOI211xp5_ASAP7_75t_R n_8257 (.A1(n_8253_o_0),
    .A2(n_8254_o_0),
    .B(n_8256_o_0),
    .C(n_7822_o_0),
    .Y(n_8257_o_0));
 AOI21xp33_ASAP7_75t_R n_8258 (.A1(n_7714_o_0),
    .A2(n_8252_o_0),
    .B(n_8257_o_0),
    .Y(n_8258_o_0));
 INVx1_ASAP7_75t_R n_8259 (.A(n_8014_o_0),
    .Y(n_8259_o_0));
 NOR2xp33_ASAP7_75t_R n_826 (.A(n_825_o_0),
    .B(n_824_o_0),
    .Y(n_826_o_0));
 INVx1_ASAP7_75t_R n_8260 (.A(n_7849_o_0),
    .Y(n_8260_o_0));
 OAI211xp5_ASAP7_75t_R n_8261 (.A1(n_7832_o_0),
    .A2(n_7821_o_0),
    .B(n_8260_o_0),
    .C(n_7837_o_0),
    .Y(n_8261_o_0));
 OAI211xp5_ASAP7_75t_R n_8262 (.A1(n_7818_o_0),
    .A2(n_7783_o_0),
    .B(n_8205_o_0),
    .C(n_7722_o_0),
    .Y(n_8262_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8263 (.A1(n_7809_o_0),
    .A2(n_8259_o_0),
    .B(n_8261_o_0),
    .C(n_8262_o_0),
    .Y(n_8263_o_0));
 NAND3xp33_ASAP7_75t_R n_8264 (.A(n_8049_o_0),
    .B(n_7991_o_0),
    .C(n_7809_o_0),
    .Y(n_8264_o_0));
 OAI311xp33_ASAP7_75t_R n_8265 (.A1(net34),
    .A2(n_7991_o_0),
    .A3(n_7796_o_0),
    .B1(n_7786_o_0),
    .C1(n_7992_o_0),
    .Y(n_8265_o_0));
 AOI31xp33_ASAP7_75t_R n_8266 (.A1(n_8264_o_0),
    .A2(n_8265_o_0),
    .A3(n_7916_o_0),
    .B(n_7910_o_0),
    .Y(n_8266_o_0));
 AOI211xp5_ASAP7_75t_R n_8267 (.A1(n_7768_o_0),
    .A2(net96),
    .B(n_7809_o_0),
    .C(n_7755_o_0),
    .Y(n_8267_o_0));
 AOI31xp33_ASAP7_75t_R n_8268 (.A1(n_7818_o_0),
    .A2(n_8171_o_0),
    .A3(n_7934_o_0),
    .B(n_8267_o_0),
    .Y(n_8268_o_0));
 OAI211xp5_ASAP7_75t_R n_8269 (.A1(n_7818_o_0),
    .A2(n_8260_o_0),
    .B(n_8268_o_0),
    .C(n_7723_o_0),
    .Y(n_8269_o_0));
 INVx3_ASAP7_75t_R n_827 (.A(ld),
    .Y(n_827_o_0));
 AOI21xp33_ASAP7_75t_R n_8270 (.A1(n_8266_o_0),
    .A2(n_8269_o_0),
    .B(n_7855_o_0),
    .Y(n_8270_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8271 (.A1(n_8263_o_0),
    .A2(n_7822_o_0),
    .B(n_8270_o_0),
    .C(n_7703_o_0),
    .Y(n_8271_o_0));
 OAI21xp33_ASAP7_75t_R n_8272 (.A1(n_7860_o_0),
    .A2(n_8258_o_0),
    .B(n_8271_o_0),
    .Y(n_8272_o_0));
 OAI21xp33_ASAP7_75t_R n_8273 (.A1(n_7906_o_0),
    .A2(n_8248_o_0),
    .B(n_8272_o_0),
    .Y(n_8273_o_0));
 XOR2xp5_ASAP7_75t_R n_8274 (.A(_01097_),
    .B(_01098_),
    .Y(n_8274_o_0));
 XNOR2xp5_ASAP7_75t_R n_8275 (.A(_01089_),
    .B(n_8274_o_0),
    .Y(n_8275_o_0));
 NOR2xp33_ASAP7_75t_R n_8276 (.A(n_3664_o_0),
    .B(n_8275_o_0),
    .Y(n_8276_o_0));
 NOR2xp33_ASAP7_75t_R n_8277 (.A(_00679_),
    .B(net),
    .Y(n_8277_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8278 (.A1(n_3664_o_0),
    .A2(n_8275_o_0),
    .B(n_8276_o_0),
    .C(net),
    .D(n_8277_o_0),
    .Y(n_8278_o_0));
 XNOR2xp5_ASAP7_75t_R n_8279 (.A(_00907_),
    .B(n_8278_o_0),
    .Y(n_8279_o_0));
 NOR2xp33_ASAP7_75t_R n_828 (.A(key[20]),
    .B(n_827_o_0),
    .Y(n_828_o_0));
 INVx1_ASAP7_75t_R n_8280 (.A(n_8279_o_0),
    .Y(n_8280_o_0));
 NAND2xp33_ASAP7_75t_R n_8281 (.A(n_3691_o_0),
    .B(n_3715_o_0),
    .Y(n_8281_o_0));
 OAI21xp33_ASAP7_75t_R n_8282 (.A1(n_3691_o_0),
    .A2(n_3715_o_0),
    .B(n_8281_o_0),
    .Y(n_8282_o_0));
 XOR2xp5_ASAP7_75t_R n_8283 (.A(_01096_),
    .B(n_8282_o_0),
    .Y(n_8283_o_0));
 NOR2xp33_ASAP7_75t_R n_8284 (.A(_00681_),
    .B(net),
    .Y(n_8284_o_0));
 INVx1_ASAP7_75t_R n_8285 (.A(n_8284_o_0),
    .Y(n_8285_o_0));
 OAI21xp33_ASAP7_75t_R n_8286 (.A1(net9),
    .A2(n_8283_o_0),
    .B(n_8285_o_0),
    .Y(n_8286_o_0));
 INVx1_ASAP7_75t_R n_8287 (.A(n_8286_o_0),
    .Y(n_8287_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8288 (.A1(net2),
    .A2(n_8283_o_0),
    .B(n_8285_o_0),
    .C(_00905_),
    .Y(n_8288_o_0));
 AOI21xp33_ASAP7_75t_R n_8289 (.A1(_00905_),
    .A2(n_8287_o_0),
    .B(n_8288_o_0),
    .Y(n_8289_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_829 (.A1(n_824_o_0),
    .A2(n_825_o_0),
    .B(n_826_o_0),
    .C(n_827_o_0),
    .D(n_828_o_0),
    .Y(n_829_o_0));
 XNOR2xp5_ASAP7_75t_R n_8290 (.A(_01097_),
    .B(n_3598_o_0),
    .Y(n_8290_o_0));
 NOR2xp33_ASAP7_75t_R n_8291 (.A(n_3606_o_0),
    .B(n_8290_o_0),
    .Y(n_8291_o_0));
 NOR2xp33_ASAP7_75t_R n_8292 (.A(_00680_),
    .B(net),
    .Y(n_8292_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8293 (.A1(n_3606_o_0),
    .A2(n_8290_o_0),
    .B(n_8291_o_0),
    .C(net),
    .D(n_8292_o_0),
    .Y(n_8293_o_0));
 NAND2xp33_ASAP7_75t_R n_8294 (.A(_00906_),
    .B(n_8293_o_0),
    .Y(n_8294_o_0));
 OAI21xp33_ASAP7_75t_R n_8295 (.A1(_00906_),
    .A2(n_8293_o_0),
    .B(n_8294_o_0),
    .Y(n_8295_o_0));
 XNOR2xp5_ASAP7_75t_R n_8296 (.A(_01007_),
    .B(_01047_),
    .Y(n_8296_o_0));
 XNOR2xp5_ASAP7_75t_R n_8297 (.A(_01093_),
    .B(_01098_),
    .Y(n_8297_o_0));
 XOR2xp5_ASAP7_75t_R n_8298 (.A(n_8296_o_0),
    .B(n_8297_o_0),
    .Y(n_8298_o_0));
 XNOR2xp5_ASAP7_75t_R n_8299 (.A(_01094_),
    .B(n_6042_o_0),
    .Y(n_8299_o_0));
 XNOR2xp5_ASAP7_75t_R n_830 (.A(_00942_),
    .B(_00974_),
    .Y(n_830_o_0));
 NOR2xp33_ASAP7_75t_R n_8300 (.A(n_8299_o_0),
    .B(n_8298_o_0),
    .Y(n_8300_o_0));
 NOR2xp33_ASAP7_75t_R n_8301 (.A(_00683_),
    .B(_00858_),
    .Y(n_8301_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8302 (.A1(n_8298_o_0),
    .A2(n_8299_o_0),
    .B(n_8300_o_0),
    .C(_00858_),
    .D(n_8301_o_0),
    .Y(n_8302_o_0));
 NAND2xp33_ASAP7_75t_R n_8303 (.A(_00903_),
    .B(n_8302_o_0),
    .Y(n_8303_o_0));
 OAI21xp5_ASAP7_75t_R n_8304 (.A1(_00903_),
    .A2(n_8302_o_0),
    .B(n_8303_o_0),
    .Y(n_8304_o_0));
 INVx1_ASAP7_75t_R n_8305 (.A(_00902_),
    .Y(n_8305_o_0));
 XNOR2xp5_ASAP7_75t_R n_8306 (.A(_01006_),
    .B(_01046_),
    .Y(n_8306_o_0));
 NAND2xp33_ASAP7_75t_R n_8307 (.A(_01093_),
    .B(n_8306_o_0),
    .Y(n_8307_o_0));
 OAI21xp33_ASAP7_75t_R n_8308 (.A1(_01093_),
    .A2(n_8306_o_0),
    .B(n_8307_o_0),
    .Y(n_8308_o_0));
 INVx1_ASAP7_75t_R n_8309 (.A(n_6018_o_0),
    .Y(n_8309_o_0));
 XNOR2xp5_ASAP7_75t_R n_831 (.A(_00910_),
    .B(n_830_o_0),
    .Y(n_831_o_0));
 OAI211xp5_ASAP7_75t_R n_8310 (.A1(_01093_),
    .A2(n_8306_o_0),
    .B(n_8307_o_0),
    .C(n_8309_o_0),
    .Y(n_8310_o_0));
 INVx1_ASAP7_75t_R n_8311 (.A(n_8310_o_0),
    .Y(n_8311_o_0));
 NOR2xp33_ASAP7_75t_R n_8312 (.A(_00584_),
    .B(_00858_),
    .Y(n_8312_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8313 (.A1(n_6018_o_0),
    .A2(n_8308_o_0),
    .B(n_8311_o_0),
    .C(net39),
    .D(n_8312_o_0),
    .Y(n_8313_o_0));
 NOR2xp33_ASAP7_75t_R n_8314 (.A(_01093_),
    .B(n_8306_o_0),
    .Y(n_8314_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8315 (.A1(_01093_),
    .A2(n_8306_o_0),
    .B(n_8314_o_0),
    .C(n_6018_o_0),
    .Y(n_8315_o_0));
 INVx1_ASAP7_75t_R n_8316 (.A(n_8312_o_0),
    .Y(n_8316_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8317 (.A1(n_8310_o_0),
    .A2(n_8315_o_0),
    .B(net3),
    .C(n_8316_o_0),
    .D(n_8305_o_0),
    .Y(n_8317_o_0));
 AOI21x1_ASAP7_75t_R n_8318 (.A1(n_8313_o_0),
    .A2(n_8305_o_0),
    .B(n_8317_o_0),
    .Y(n_8318_o_0));
 XNOR2xp5_ASAP7_75t_R n_8319 (.A(_01091_),
    .B(_01098_),
    .Y(n_8319_o_0));
 XNOR2xp5_ASAP7_75t_R n_832 (.A(_00417_),
    .B(_00878_),
    .Y(n_832_o_0));
 XNOR2xp5_ASAP7_75t_R n_8320 (.A(_01044_),
    .B(_01090_),
    .Y(n_8320_o_0));
 NAND2xp33_ASAP7_75t_R n_8321 (.A(n_3653_o_0),
    .B(n_8320_o_0),
    .Y(n_8321_o_0));
 OAI21xp33_ASAP7_75t_R n_8322 (.A1(n_8320_o_0),
    .A2(n_3653_o_0),
    .B(n_8321_o_0),
    .Y(n_8322_o_0));
 XOR2xp5_ASAP7_75t_R n_8323 (.A(_01091_),
    .B(_01098_),
    .Y(n_8323_o_0));
 OAI211xp5_ASAP7_75t_R n_8324 (.A1(n_8320_o_0),
    .A2(n_3653_o_0),
    .B(n_8321_o_0),
    .C(n_8323_o_0),
    .Y(n_8324_o_0));
 INVx1_ASAP7_75t_R n_8325 (.A(n_8324_o_0),
    .Y(n_8325_o_0));
 NOR2xp33_ASAP7_75t_R n_8326 (.A(_00582_),
    .B(net39),
    .Y(n_8326_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8327 (.A1(n_8319_o_0),
    .A2(n_8322_o_0),
    .B(n_8325_o_0),
    .C(net39),
    .D(n_8326_o_0),
    .Y(n_8327_o_0));
 NOR2xp33_ASAP7_75t_R n_8328 (.A(n_3653_o_0),
    .B(n_8320_o_0),
    .Y(n_8328_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8329 (.A1(n_8320_o_0),
    .A2(n_3653_o_0),
    .B(n_8328_o_0),
    .C(n_8319_o_0),
    .Y(n_8329_o_0));
 INVx1_ASAP7_75t_R n_833 (.A(n_832_o_0),
    .Y(n_833_o_0));
 INVx1_ASAP7_75t_R n_8330 (.A(n_8326_o_0),
    .Y(n_8330_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8331 (.A1(n_8324_o_0),
    .A2(n_8329_o_0),
    .B(net3),
    .C(n_8330_o_0),
    .D(_00900_),
    .Y(n_8331_o_0));
 AOI21x1_ASAP7_75t_R n_8332 (.A1(_00900_),
    .A2(n_8327_o_0),
    .B(n_8331_o_0),
    .Y(n_8332_o_0));
 NAND2xp33_ASAP7_75t_R n_8333 (.A(n_6004_o_0),
    .B(n_8323_o_0),
    .Y(n_8333_o_0));
 OAI21xp33_ASAP7_75t_R n_8334 (.A1(n_6004_o_0),
    .A2(n_8323_o_0),
    .B(n_8333_o_0),
    .Y(n_8334_o_0));
 NAND2xp33_ASAP7_75t_R n_8335 (.A(_01092_),
    .B(n_3629_o_0),
    .Y(n_8335_o_0));
 OAI21xp33_ASAP7_75t_R n_8336 (.A1(_01092_),
    .A2(n_3629_o_0),
    .B(n_8335_o_0),
    .Y(n_8336_o_0));
 OAI21xp33_ASAP7_75t_R n_8337 (.A1(n_8336_o_0),
    .A2(n_8334_o_0),
    .B(net39),
    .Y(n_8337_o_0));
 AOI21xp33_ASAP7_75t_R n_8338 (.A1(n_8334_o_0),
    .A2(n_8336_o_0),
    .B(n_8337_o_0),
    .Y(n_8338_o_0));
 NOR2xp33_ASAP7_75t_R n_8339 (.A(n_6004_o_0),
    .B(n_8323_o_0),
    .Y(n_8339_o_0));
 AO21x1_ASAP7_75t_R n_834 (.A1(n_831_o_0),
    .A2(n_833_o_0),
    .B(ld),
    .Y(n_834_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8340 (.A1(n_6004_o_0),
    .A2(n_8323_o_0),
    .B(n_8339_o_0),
    .C(n_8336_o_0),
    .Y(n_8340_o_0));
 XNOR2xp5_ASAP7_75t_R n_8341 (.A(n_8319_o_0),
    .B(n_6004_o_0),
    .Y(n_8341_o_0));
 XOR2xp5_ASAP7_75t_R n_8342 (.A(_01092_),
    .B(n_3629_o_0),
    .Y(n_8342_o_0));
 AOI21xp33_ASAP7_75t_R n_8343 (.A1(n_8341_o_0),
    .A2(n_8342_o_0),
    .B(net5),
    .Y(n_8343_o_0));
 AOI221xp5_ASAP7_75t_R n_8344 (.A1(net1),
    .A2(_00581_),
    .B1(n_8340_o_0),
    .B2(n_8343_o_0),
    .C(_00901_),
    .Y(n_8344_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8345 (.A1(net5),
    .A2(_00581_),
    .B(n_8338_o_0),
    .C(_00901_),
    .D(n_8344_o_0),
    .Y(n_8345_o_0));
 NOR2xp33_ASAP7_75t_R n_8346 (.A(n_8332_o_0),
    .B(n_8345_o_0),
    .Y(n_8346_o_0));
 NOR2xp33_ASAP7_75t_R n_8347 (.A(n_8318_o_0),
    .B(n_8346_o_0),
    .Y(n_8347_o_0));
 NAND2xp33_ASAP7_75t_R n_8348 (.A(n_8318_o_0),
    .B(n_8346_o_0),
    .Y(n_8348_o_0));
 INVx1_ASAP7_75t_R n_8349 (.A(n_8348_o_0),
    .Y(n_8349_o_0));
 NOR3xp33_ASAP7_75t_R n_835 (.A(n_831_o_0),
    .B(n_833_o_0),
    .C(ld),
    .Y(n_835_o_0));
 INVx1_ASAP7_75t_R n_8350 (.A(_01094_),
    .Y(n_8350_o_0));
 NOR2xp33_ASAP7_75t_R n_8351 (.A(n_8350_o_0),
    .B(n_6042_o_0),
    .Y(n_8351_o_0));
 XNOR2xp5_ASAP7_75t_R n_8352 (.A(n_8296_o_0),
    .B(n_8297_o_0),
    .Y(n_8352_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8353 (.A1(n_6042_o_0),
    .A2(n_8350_o_0),
    .B(n_8351_o_0),
    .C(n_8352_o_0),
    .Y(n_8353_o_0));
 NAND2xp33_ASAP7_75t_R n_8354 (.A(n_8299_o_0),
    .B(n_8298_o_0),
    .Y(n_8354_o_0));
 INVx1_ASAP7_75t_R n_8355 (.A(n_8301_o_0),
    .Y(n_8355_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8356 (.A1(n_8353_o_0),
    .A2(n_8354_o_0),
    .B(net3),
    .C(n_8355_o_0),
    .D(n_1393_o_0),
    .Y(n_8356_o_0));
 AOI21x1_ASAP7_75t_R n_8357 (.A1(n_1393_o_0),
    .A2(n_8302_o_0),
    .B(n_8356_o_0),
    .Y(n_8357_o_0));
 INVx2_ASAP7_75t_R n_8358 (.A(n_8357_o_0),
    .Y(n_8358_o_0));
 INVx1_ASAP7_75t_R n_8359 (.A(_00581_),
    .Y(n_8359_o_0));
 O2A1O1Ixp5_ASAP7_75t_R n_836 (.A1(n_827_o_0),
    .A2(key[18]),
    .B(n_834_o_0),
    .C(n_835_o_0),
    .Y(n_836_o_0));
 NOR2xp33_ASAP7_75t_R n_8360 (.A(n_8341_o_0),
    .B(n_8342_o_0),
    .Y(n_8360_o_0));
 INVx1_ASAP7_75t_R n_8361 (.A(_00901_),
    .Y(n_8361_o_0));
 OAI221xp5_ASAP7_75t_R n_8362 (.A1(net39),
    .A2(n_8359_o_0),
    .B1(n_8337_o_0),
    .B2(n_8360_o_0),
    .C(n_8361_o_0),
    .Y(n_8362_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8363 (.A1(net2),
    .A2(_00581_),
    .B(n_8338_o_0),
    .C(_00901_),
    .Y(n_8363_o_0));
 AOI21xp33_ASAP7_75t_R n_8364 (.A1(n_8362_o_0),
    .A2(n_8363_o_0),
    .B(n_8332_o_0),
    .Y(n_8364_o_0));
 AO21x1_ASAP7_75t_R n_8365 (.A1(n_8313_o_0),
    .A2(n_8305_o_0),
    .B(n_8317_o_0),
    .Y(n_8365_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8366 (.A1(n_8332_o_0),
    .A2(n_8345_o_0),
    .B(n_8364_o_0),
    .C(n_8365_o_0),
    .Y(n_8366_o_0));
 NAND2xp33_ASAP7_75t_R n_8367 (.A(n_8358_o_0),
    .B(n_8366_o_0),
    .Y(n_8367_o_0));
 OAI211xp5_ASAP7_75t_R n_8368 (.A1(n_8334_o_0),
    .A2(n_8336_o_0),
    .B(n_8340_o_0),
    .C(net39),
    .Y(n_8368_o_0));
 NAND2xp33_ASAP7_75t_R n_8369 (.A(_00581_),
    .B(n_3021_o_0),
    .Y(n_8369_o_0));
 XNOR2xp5_ASAP7_75t_R n_837 (.A(_00940_),
    .B(_00972_),
    .Y(n_837_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8370 (.A1(n_8368_o_0),
    .A2(n_8369_o_0),
    .B(n_8361_o_0),
    .C(n_8362_o_0),
    .Y(n_8370_o_0));
 NAND2xp33_ASAP7_75t_R n_8371 (.A(n_8332_o_0),
    .B(n_8370_o_0),
    .Y(n_8371_o_0));
 NAND3xp33_ASAP7_75t_R n_8372 (.A(n_8304_o_0),
    .B(n_8371_o_0),
    .C(net73),
    .Y(n_8372_o_0));
 OAI21xp33_ASAP7_75t_R n_8373 (.A1(n_8349_o_0),
    .A2(n_8367_o_0),
    .B(n_8372_o_0),
    .Y(n_8373_o_0));
 XOR2xp5_ASAP7_75t_R n_8374 (.A(_01094_),
    .B(_01098_),
    .Y(n_8374_o_0));
 XNOR2xp5_ASAP7_75t_R n_8375 (.A(n_3597_o_0),
    .B(n_8374_o_0),
    .Y(n_8375_o_0));
 XNOR2xp5_ASAP7_75t_R n_8376 (.A(_01095_),
    .B(n_5996_o_0),
    .Y(n_8376_o_0));
 NOR2xp33_ASAP7_75t_R n_8377 (.A(n_8376_o_0),
    .B(n_8375_o_0),
    .Y(n_8377_o_0));
 NOR2xp33_ASAP7_75t_R n_8378 (.A(_00682_),
    .B(net39),
    .Y(n_8378_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8379 (.A1(n_8375_o_0),
    .A2(n_8376_o_0),
    .B(n_8377_o_0),
    .C(net39),
    .D(n_8378_o_0),
    .Y(n_8379_o_0));
 XOR2xp5_ASAP7_75t_R n_838 (.A(_00439_),
    .B(_00876_),
    .Y(n_838_o_0));
 XOR2x1_ASAP7_75t_R n_8380 (.A(_00904_),
    .Y(n_8380_o_0),
    .B(n_8379_o_0));
 INVx1_ASAP7_75t_R n_8381 (.A(n_8380_o_0),
    .Y(n_8381_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8382 (.A1(n_8304_o_0),
    .A2(n_8347_o_0),
    .B(n_8373_o_0),
    .C(n_8381_o_0),
    .Y(n_8382_o_0));
 NOR2xp33_ASAP7_75t_R n_8383 (.A(net38),
    .B(n_8365_o_0),
    .Y(n_8383_o_0));
 AO21x1_ASAP7_75t_R n_8384 (.A1(n_8327_o_0),
    .A2(_00900_),
    .B(n_8331_o_0),
    .Y(n_8384_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8385 (.A1(_00900_),
    .A2(n_8327_o_0),
    .B(n_8331_o_0),
    .C(n_8370_o_0),
    .Y(n_8385_o_0));
 OAI21xp33_ASAP7_75t_R n_8386 (.A1(n_8384_o_0),
    .A2(n_8370_o_0),
    .B(n_8385_o_0),
    .Y(n_8386_o_0));
 OAI21xp33_ASAP7_75t_R n_8387 (.A1(n_8318_o_0),
    .A2(n_8386_o_0),
    .B(n_8304_o_0),
    .Y(n_8387_o_0));
 NAND2xp33_ASAP7_75t_R n_8388 (.A(n_8369_o_0),
    .B(n_8368_o_0),
    .Y(n_8388_o_0));
 OAI211xp5_ASAP7_75t_R n_8389 (.A1(_00901_),
    .A2(n_8388_o_0),
    .B(n_8332_o_0),
    .C(n_8363_o_0),
    .Y(n_8389_o_0));
 INVx1_ASAP7_75t_R n_839 (.A(_00908_),
    .Y(n_839_o_0));
 AOI21xp33_ASAP7_75t_R n_8390 (.A1(n_8385_o_0),
    .A2(n_8389_o_0),
    .B(n_8365_o_0),
    .Y(n_8390_o_0));
 INVx1_ASAP7_75t_R n_8391 (.A(n_8390_o_0),
    .Y(n_8391_o_0));
 NAND2xp33_ASAP7_75t_R n_8392 (.A(_00904_),
    .B(n_8379_o_0),
    .Y(n_8392_o_0));
 OAI21xp33_ASAP7_75t_R n_8393 (.A1(_00904_),
    .A2(n_8379_o_0),
    .B(n_8392_o_0),
    .Y(n_8393_o_0));
 AOI21xp33_ASAP7_75t_R n_8394 (.A1(n_8358_o_0),
    .A2(n_8391_o_0),
    .B(n_8393_o_0),
    .Y(n_8394_o_0));
 OAI21xp33_ASAP7_75t_R n_8395 (.A1(n_8383_o_0),
    .A2(n_8387_o_0),
    .B(n_8394_o_0),
    .Y(n_8395_o_0));
 NAND2xp33_ASAP7_75t_R n_8396 (.A(n_8318_o_0),
    .B(n_8384_o_0),
    .Y(n_8396_o_0));
 INVx1_ASAP7_75t_R n_8397 (.A(n_8396_o_0),
    .Y(n_8397_o_0));
 AOI21xp33_ASAP7_75t_R n_8398 (.A1(n_8332_o_0),
    .A2(n_8345_o_0),
    .B(n_8318_o_0),
    .Y(n_8398_o_0));
 NAND2xp33_ASAP7_75t_R n_8399 (.A(n_8345_o_0),
    .B(n_8384_o_0),
    .Y(n_8399_o_0));
 NAND2xp33_ASAP7_75t_R n_840 (.A(n_839_o_0),
    .B(n_838_o_0),
    .Y(n_840_o_0));
 NOR2xp33_ASAP7_75t_R n_8400 (.A(n_8318_o_0),
    .B(n_8345_o_0),
    .Y(n_8400_o_0));
 INVx1_ASAP7_75t_R n_8401 (.A(n_8400_o_0),
    .Y(n_8401_o_0));
 OAI211xp5_ASAP7_75t_R n_8402 (.A1(n_8365_o_0),
    .A2(n_8399_o_0),
    .B(n_8401_o_0),
    .C(n_8304_o_0),
    .Y(n_8402_o_0));
 OAI31xp33_ASAP7_75t_R n_8403 (.A1(n_8357_o_0),
    .A2(n_8397_o_0),
    .A3(n_8398_o_0),
    .B(n_8402_o_0),
    .Y(n_8403_o_0));
 OAI211xp5_ASAP7_75t_R n_8404 (.A1(n_8384_o_0),
    .A2(n_8318_o_0),
    .B(net66),
    .C(n_8357_o_0),
    .Y(n_8404_o_0));
 NAND2xp33_ASAP7_75t_R n_8405 (.A(n_8332_o_0),
    .B(n_8345_o_0),
    .Y(n_8405_o_0));
 NAND2xp33_ASAP7_75t_R n_8406 (.A(n_8318_o_0),
    .B(n_8384_o_0),
    .Y(n_8406_o_0));
 NOR2xp33_ASAP7_75t_R n_8407 (.A(_00903_),
    .B(n_8302_o_0),
    .Y(n_8407_o_0));
 AOI21xp5_ASAP7_75t_R n_8408 (.A1(_00903_),
    .A2(n_8302_o_0),
    .B(n_8407_o_0),
    .Y(n_8408_o_0));
 OAI211xp5_ASAP7_75t_R n_8409 (.A1(n_8405_o_0),
    .A2(n_8318_o_0),
    .B(n_8406_o_0),
    .C(n_8408_o_0),
    .Y(n_8409_o_0));
 OAI21xp33_ASAP7_75t_R n_841 (.A1(n_838_o_0),
    .A2(n_839_o_0),
    .B(n_840_o_0),
    .Y(n_841_o_0));
 AOI21xp33_ASAP7_75t_R n_8410 (.A1(n_8404_o_0),
    .A2(n_8409_o_0),
    .B(n_8380_o_0),
    .Y(n_8410_o_0));
 AOI211xp5_ASAP7_75t_R n_8411 (.A1(n_8403_o_0),
    .A2(n_8380_o_0),
    .B(n_8295_o_0),
    .C(n_8410_o_0),
    .Y(n_8411_o_0));
 AOI31xp33_ASAP7_75t_R n_8412 (.A1(n_8295_o_0),
    .A2(n_8382_o_0),
    .A3(n_8395_o_0),
    .B(n_8411_o_0),
    .Y(n_8412_o_0));
 XNOR2xp5_ASAP7_75t_R n_8413 (.A(_00906_),
    .B(n_8293_o_0),
    .Y(n_8413_o_0));
 INVx1_ASAP7_75t_R n_8414 (.A(n_8413_o_0),
    .Y(n_8414_o_0));
 AND2x2_ASAP7_75t_R n_8415 (.A(_00903_),
    .B(n_8302_o_0),
    .Y(n_8415_o_0));
 OAI22xp33_ASAP7_75t_R n_8416 (.A1(n_8415_o_0),
    .A2(n_8407_o_0),
    .B1(n_8384_o_0),
    .B2(n_8318_o_0),
    .Y(n_8416_o_0));
 AOI21xp33_ASAP7_75t_R n_8417 (.A1(n_8384_o_0),
    .A2(net38),
    .B(n_8416_o_0),
    .Y(n_8417_o_0));
 NAND2xp33_ASAP7_75t_R n_8418 (.A(n_8370_o_0),
    .B(n_8384_o_0),
    .Y(n_8418_o_0));
 NAND2xp33_ASAP7_75t_R n_8419 (.A(n_8332_o_0),
    .B(n_8365_o_0),
    .Y(n_8419_o_0));
 NAND2xp33_ASAP7_75t_R n_842 (.A(n_837_o_0),
    .B(n_841_o_0),
    .Y(n_842_o_0));
 AOI21xp33_ASAP7_75t_R n_8420 (.A1(n_8418_o_0),
    .A2(n_8419_o_0),
    .B(n_8304_o_0),
    .Y(n_8420_o_0));
 NOR2xp33_ASAP7_75t_R n_8421 (.A(n_8365_o_0),
    .B(n_8405_o_0),
    .Y(n_8421_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8422 (.A1(n_8389_o_0),
    .A2(n_8385_o_0),
    .B(n_8318_o_0),
    .C(n_8357_o_0),
    .Y(n_8422_o_0));
 OAI21xp33_ASAP7_75t_R n_8423 (.A1(n_8318_o_0),
    .A2(n_8371_o_0),
    .B(n_8358_o_0),
    .Y(n_8423_o_0));
 OAI221xp5_ASAP7_75t_R n_8424 (.A1(n_8421_o_0),
    .A2(n_8422_o_0),
    .B1(n_8423_o_0),
    .B2(n_8349_o_0),
    .C(n_8393_o_0),
    .Y(n_8424_o_0));
 OAI31xp33_ASAP7_75t_R n_8425 (.A1(n_8381_o_0),
    .A2(n_8417_o_0),
    .A3(n_8420_o_0),
    .B(n_8424_o_0),
    .Y(n_8425_o_0));
 INVx1_ASAP7_75t_R n_8426 (.A(n_8295_o_0),
    .Y(n_8426_o_0));
 AOI21xp33_ASAP7_75t_R n_8427 (.A1(n_8332_o_0),
    .A2(n_8345_o_0),
    .B(n_8365_o_0),
    .Y(n_8427_o_0));
 NOR3xp33_ASAP7_75t_R n_8428 (.A(n_8365_o_0),
    .B(net66),
    .C(n_8332_o_0),
    .Y(n_8428_o_0));
 INVx1_ASAP7_75t_R n_8429 (.A(n_8428_o_0),
    .Y(n_8429_o_0));
 INVx1_ASAP7_75t_R n_843 (.A(n_837_o_0),
    .Y(n_843_o_0));
 NOR2xp33_ASAP7_75t_R n_8430 (.A(n_8332_o_0),
    .B(n_8318_o_0),
    .Y(n_8430_o_0));
 INVx1_ASAP7_75t_R n_8431 (.A(n_8430_o_0),
    .Y(n_8431_o_0));
 AOI31xp33_ASAP7_75t_R n_8432 (.A1(n_8304_o_0),
    .A2(n_8429_o_0),
    .A3(n_8431_o_0),
    .B(n_8393_o_0),
    .Y(n_8432_o_0));
 OAI21xp33_ASAP7_75t_R n_8433 (.A1(n_8427_o_0),
    .A2(n_8367_o_0),
    .B(n_8432_o_0),
    .Y(n_8433_o_0));
 NOR2xp67_ASAP7_75t_R n_8434 (.A(n_8332_o_0),
    .B(n_8370_o_0),
    .Y(n_8434_o_0));
 OAI21xp33_ASAP7_75t_R n_8435 (.A1(n_8318_o_0),
    .A2(n_8434_o_0),
    .B(n_8408_o_0),
    .Y(n_8435_o_0));
 NAND2xp33_ASAP7_75t_R n_8436 (.A(n_8304_o_0),
    .B(n_8396_o_0),
    .Y(n_8436_o_0));
 OAI211xp5_ASAP7_75t_R n_8437 (.A1(n_8435_o_0),
    .A2(n_8428_o_0),
    .B(n_8436_o_0),
    .C(n_8381_o_0),
    .Y(n_8437_o_0));
 NAND2xp33_ASAP7_75t_R n_8438 (.A(_01096_),
    .B(n_8282_o_0),
    .Y(n_8438_o_0));
 OAI21xp33_ASAP7_75t_R n_8439 (.A1(_01096_),
    .A2(n_8282_o_0),
    .B(n_8438_o_0),
    .Y(n_8439_o_0));
 OAI211xp5_ASAP7_75t_R n_844 (.A1(n_838_o_0),
    .A2(n_839_o_0),
    .B(n_840_o_0),
    .C(n_843_o_0),
    .Y(n_844_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8440 (.A1(n_8439_o_0),
    .A2(net),
    .B(n_8284_o_0),
    .C(_00905_),
    .Y(n_8440_o_0));
 OAI21xp33_ASAP7_75t_R n_8441 (.A1(_00905_),
    .A2(n_8286_o_0),
    .B(n_8440_o_0),
    .Y(n_8441_o_0));
 INVx1_ASAP7_75t_R n_8442 (.A(n_8441_o_0),
    .Y(n_8442_o_0));
 AOI31xp33_ASAP7_75t_R n_8443 (.A1(n_8426_o_0),
    .A2(n_8433_o_0),
    .A3(n_8437_o_0),
    .B(n_8442_o_0),
    .Y(n_8443_o_0));
 OAI21xp33_ASAP7_75t_R n_8444 (.A1(n_8414_o_0),
    .A2(n_8425_o_0),
    .B(n_8443_o_0),
    .Y(n_8444_o_0));
 OAI21xp33_ASAP7_75t_R n_8445 (.A1(n_8289_o_0),
    .A2(n_8412_o_0),
    .B(n_8444_o_0),
    .Y(n_8445_o_0));
 INVx1_ASAP7_75t_R n_8446 (.A(n_8289_o_0),
    .Y(n_8446_o_0));
 NAND2xp33_ASAP7_75t_R n_8447 (.A(n_8332_o_0),
    .B(n_8318_o_0),
    .Y(n_8447_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8448 (.A1(net73),
    .A2(n_8346_o_0),
    .B(n_8447_o_0),
    .C(n_8304_o_0),
    .Y(n_8448_o_0));
 OAI21xp33_ASAP7_75t_R n_8449 (.A1(n_8358_o_0),
    .A2(n_8348_o_0),
    .B(n_8393_o_0),
    .Y(n_8449_o_0));
 NAND2xp33_ASAP7_75t_R n_845 (.A(key[16]),
    .B(ld),
    .Y(n_845_o_0));
 NOR2xp33_ASAP7_75t_R n_8450 (.A(n_8365_o_0),
    .B(n_8434_o_0),
    .Y(n_8450_o_0));
 OAI21xp33_ASAP7_75t_R n_8451 (.A1(n_8318_o_0),
    .A2(n_8399_o_0),
    .B(n_8304_o_0),
    .Y(n_8451_o_0));
 NOR2xp33_ASAP7_75t_R n_8452 (.A(n_8450_o_0),
    .B(n_8451_o_0),
    .Y(n_8452_o_0));
 NOR2xp33_ASAP7_75t_R n_8453 (.A(n_8318_o_0),
    .B(net66),
    .Y(n_8453_o_0));
 INVx1_ASAP7_75t_R n_8454 (.A(n_8453_o_0),
    .Y(n_8454_o_0));
 INVx1_ASAP7_75t_R n_8455 (.A(n_8386_o_0),
    .Y(n_8455_o_0));
 AOI21xp33_ASAP7_75t_R n_8456 (.A1(n_8318_o_0),
    .A2(n_8455_o_0),
    .B(n_8408_o_0),
    .Y(n_8456_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8457 (.A1(n_8358_o_0),
    .A2(n_8454_o_0),
    .B(n_8456_o_0),
    .C(n_8380_o_0),
    .Y(n_8457_o_0));
 OAI31xp33_ASAP7_75t_R n_8458 (.A1(n_8448_o_0),
    .A2(n_8449_o_0),
    .A3(n_8452_o_0),
    .B(n_8457_o_0),
    .Y(n_8458_o_0));
 NAND3xp33_ASAP7_75t_R n_8459 (.A(n_8399_o_0),
    .B(n_8365_o_0),
    .C(n_8304_o_0),
    .Y(n_8459_o_0));
 INVx1_ASAP7_75t_R n_846 (.A(n_845_o_0),
    .Y(n_846_o_0));
 NAND3xp33_ASAP7_75t_R n_8460 (.A(n_8346_o_0),
    .B(n_8358_o_0),
    .C(n_8365_o_0),
    .Y(n_8460_o_0));
 INVx1_ASAP7_75t_R n_8461 (.A(n_8393_o_0),
    .Y(n_8461_o_0));
 NAND4xp25_ASAP7_75t_R n_8462 (.A(n_8459_o_0),
    .B(n_8460_o_0),
    .C(n_8372_o_0),
    .D(n_8461_o_0),
    .Y(n_8462_o_0));
 NOR2xp33_ASAP7_75t_R n_8463 (.A(n_8318_o_0),
    .B(n_8399_o_0),
    .Y(n_8463_o_0));
 AOI21xp33_ASAP7_75t_R n_8464 (.A1(n_8332_o_0),
    .A2(n_8370_o_0),
    .B(n_8365_o_0),
    .Y(n_8464_o_0));
 OAI31xp33_ASAP7_75t_R n_8465 (.A1(n_8357_o_0),
    .A2(n_8463_o_0),
    .A3(n_8464_o_0),
    .B(n_8381_o_0),
    .Y(n_8465_o_0));
 NAND3xp33_ASAP7_75t_R n_8466 (.A(n_8346_o_0),
    .B(n_8365_o_0),
    .C(n_8357_o_0),
    .Y(n_8466_o_0));
 NAND2xp33_ASAP7_75t_R n_8467 (.A(n_8441_o_0),
    .B(n_8466_o_0),
    .Y(n_8467_o_0));
 OAI22xp33_ASAP7_75t_R n_8468 (.A1(n_8462_o_0),
    .A2(n_8446_o_0),
    .B1(n_8465_o_0),
    .B2(n_8467_o_0),
    .Y(n_8468_o_0));
 AOI21xp33_ASAP7_75t_R n_8469 (.A1(n_8446_o_0),
    .A2(n_8458_o_0),
    .B(n_8468_o_0),
    .Y(n_8469_o_0));
 AOI31xp67_ASAP7_75t_R n_847 (.A1(n_827_o_0),
    .A2(n_842_o_0),
    .A3(n_844_o_0),
    .B(n_846_o_0),
    .Y(n_847_o_0));
 NAND3xp33_ASAP7_75t_R n_8470 (.A(net66),
    .B(n_8318_o_0),
    .C(n_8332_o_0),
    .Y(n_8470_o_0));
 NAND2xp33_ASAP7_75t_R n_8471 (.A(n_8441_o_0),
    .B(n_8393_o_0),
    .Y(n_8471_o_0));
 AOI31xp33_ASAP7_75t_R n_8472 (.A1(n_8358_o_0),
    .A2(n_8431_o_0),
    .A3(n_8470_o_0),
    .B(n_8471_o_0),
    .Y(n_8472_o_0));
 NOR2xp33_ASAP7_75t_R n_8473 (.A(n_8318_o_0),
    .B(n_8370_o_0),
    .Y(n_8473_o_0));
 INVx1_ASAP7_75t_R n_8474 (.A(n_8473_o_0),
    .Y(n_8474_o_0));
 NAND2xp33_ASAP7_75t_R n_8475 (.A(n_8474_o_0),
    .B(n_8456_o_0),
    .Y(n_8475_o_0));
 NAND3xp33_ASAP7_75t_R n_8476 (.A(n_8365_o_0),
    .B(net66),
    .C(n_8332_o_0),
    .Y(n_8476_o_0));
 INVx1_ASAP7_75t_R n_8477 (.A(n_8476_o_0),
    .Y(n_8477_o_0));
 AOI21xp33_ASAP7_75t_R n_8478 (.A1(n_8365_o_0),
    .A2(n_8386_o_0),
    .B(n_8304_o_0),
    .Y(n_8478_o_0));
 AO21x1_ASAP7_75t_R n_8479 (.A1(n_8357_o_0),
    .A2(n_8477_o_0),
    .B(n_8478_o_0),
    .Y(n_8479_o_0));
 XNOR2xp5_ASAP7_75t_R n_848 (.A(_00941_),
    .B(_00973_),
    .Y(n_848_o_0));
 NAND3xp33_ASAP7_75t_R n_8480 (.A(n_8434_o_0),
    .B(n_8357_o_0),
    .C(net73),
    .Y(n_8480_o_0));
 INVx1_ASAP7_75t_R n_8481 (.A(n_8480_o_0),
    .Y(n_8481_o_0));
 OAI21xp33_ASAP7_75t_R n_8482 (.A1(n_8380_o_0),
    .A2(n_8409_o_0),
    .B(n_8446_o_0),
    .Y(n_8482_o_0));
 AOI211xp5_ASAP7_75t_R n_8483 (.A1(n_8479_o_0),
    .A2(n_8461_o_0),
    .B(n_8481_o_0),
    .C(n_8482_o_0),
    .Y(n_8483_o_0));
 NAND2xp33_ASAP7_75t_R n_8484 (.A(n_8370_o_0),
    .B(n_8384_o_0),
    .Y(n_8484_o_0));
 NAND2xp33_ASAP7_75t_R n_8485 (.A(n_8318_o_0),
    .B(n_8484_o_0),
    .Y(n_8485_o_0));
 AOI21xp33_ASAP7_75t_R n_8486 (.A1(n_8466_o_0),
    .A2(n_8485_o_0),
    .B(n_8358_o_0),
    .Y(n_8486_o_0));
 AOI21xp33_ASAP7_75t_R n_8487 (.A1(n_8365_o_0),
    .A2(n_8399_o_0),
    .B(n_8304_o_0),
    .Y(n_8487_o_0));
 NOR4xp25_ASAP7_75t_R n_8488 (.A(n_8486_o_0),
    .B(n_8487_o_0),
    .C(n_8442_o_0),
    .D(n_8381_o_0),
    .Y(n_8488_o_0));
 AOI211xp5_ASAP7_75t_R n_8489 (.A1(n_8472_o_0),
    .A2(n_8475_o_0),
    .B(n_8483_o_0),
    .C(n_8488_o_0),
    .Y(n_8489_o_0));
 INVx1_ASAP7_75t_R n_849 (.A(n_848_o_0),
    .Y(n_849_o_0));
 OAI221xp5_ASAP7_75t_R n_8490 (.A1(n_8426_o_0),
    .A2(n_8469_o_0),
    .B1(n_8489_o_0),
    .B2(n_8413_o_0),
    .C(n_8280_o_0),
    .Y(n_8490_o_0));
 OAI21xp33_ASAP7_75t_R n_8491 (.A1(n_8280_o_0),
    .A2(n_8445_o_0),
    .B(n_8490_o_0),
    .Y(n_8491_o_0));
 INVx1_ASAP7_75t_R n_8492 (.A(n_8398_o_0),
    .Y(n_8492_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8493 (.A1(n_8389_o_0),
    .A2(n_8385_o_0),
    .B(n_8365_o_0),
    .C(n_8492_o_0),
    .Y(n_8493_o_0));
 OAI22xp33_ASAP7_75t_R n_8494 (.A1(n_8493_o_0),
    .A2(n_8357_o_0),
    .B1(n_8450_o_0),
    .B2(n_8451_o_0),
    .Y(n_8494_o_0));
 OAI21xp33_ASAP7_75t_R n_8495 (.A1(net45),
    .A2(n_8318_o_0),
    .B(n_8357_o_0),
    .Y(n_8495_o_0));
 INVx1_ASAP7_75t_R n_8496 (.A(n_8495_o_0),
    .Y(n_8496_o_0));
 AOI311xp33_ASAP7_75t_R n_8497 (.A1(n_8408_o_0),
    .A2(net45),
    .A3(net73),
    .B(n_8381_o_0),
    .C(n_8496_o_0),
    .Y(n_8497_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8498 (.A1(n_8381_o_0),
    .A2(n_8481_o_0),
    .B(n_8494_o_0),
    .C(n_8497_o_0),
    .Y(n_8498_o_0));
 AOI211xp5_ASAP7_75t_R n_8499 (.A1(n_8365_o_0),
    .A2(net45),
    .B(n_8408_o_0),
    .C(net67),
    .Y(n_8499_o_0));
 XOR2xp5_ASAP7_75t_R n_850 (.A(_00440_),
    .B(_00877_),
    .Y(n_850_o_0));
 AOI31xp33_ASAP7_75t_R n_8500 (.A1(n_8358_o_0),
    .A2(n_8366_o_0),
    .A3(n_8429_o_0),
    .B(n_8499_o_0),
    .Y(n_8500_o_0));
 NAND2xp33_ASAP7_75t_R n_8501 (.A(n_8332_o_0),
    .B(n_8345_o_0),
    .Y(n_8501_o_0));
 AOI21xp33_ASAP7_75t_R n_8502 (.A1(n_8386_o_0),
    .A2(net73),
    .B(n_8416_o_0),
    .Y(n_8502_o_0));
 AOI31xp33_ASAP7_75t_R n_8503 (.A1(n_8358_o_0),
    .A2(n_8431_o_0),
    .A3(n_8501_o_0),
    .B(n_8502_o_0),
    .Y(n_8503_o_0));
 OAI221xp5_ASAP7_75t_R n_8504 (.A1(n_8381_o_0),
    .A2(n_8500_o_0),
    .B1(n_8461_o_0),
    .B2(n_8503_o_0),
    .C(n_8426_o_0),
    .Y(n_8504_o_0));
 OAI21xp33_ASAP7_75t_R n_8505 (.A1(n_8426_o_0),
    .A2(n_8498_o_0),
    .B(n_8504_o_0),
    .Y(n_8505_o_0));
 NAND2xp33_ASAP7_75t_R n_8506 (.A(n_8318_o_0),
    .B(n_8358_o_0),
    .Y(n_8506_o_0));
 NAND3xp33_ASAP7_75t_R n_8507 (.A(n_8474_o_0),
    .B(n_8418_o_0),
    .C(n_8304_o_0),
    .Y(n_8507_o_0));
 OAI21xp33_ASAP7_75t_R n_8508 (.A1(n_8434_o_0),
    .A2(n_8506_o_0),
    .B(n_8507_o_0),
    .Y(n_8508_o_0));
 INVx1_ASAP7_75t_R n_8509 (.A(n_8508_o_0),
    .Y(n_8509_o_0));
 XNOR2xp5_ASAP7_75t_R n_851 (.A(_00909_),
    .B(n_850_o_0),
    .Y(n_851_o_0));
 OAI21xp33_ASAP7_75t_R n_8510 (.A1(n_8318_o_0),
    .A2(n_8434_o_0),
    .B(n_8357_o_0),
    .Y(n_8510_o_0));
 INVx1_ASAP7_75t_R n_8511 (.A(n_8510_o_0),
    .Y(n_8511_o_0));
 NAND2xp33_ASAP7_75t_R n_8512 (.A(net67),
    .B(n_8318_o_0),
    .Y(n_8512_o_0));
 AO21x1_ASAP7_75t_R n_8513 (.A1(n_8478_o_0),
    .A2(n_8406_o_0),
    .B(n_8381_o_0),
    .Y(n_8513_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8514 (.A1(n_8511_o_0),
    .A2(n_8512_o_0),
    .B(n_8513_o_0),
    .C(n_8295_o_0),
    .Y(n_8514_o_0));
 AOI211xp5_ASAP7_75t_R n_8515 (.A1(n_8381_o_0),
    .A2(n_8509_o_0),
    .B(n_8514_o_0),
    .C(n_8442_o_0),
    .Y(n_8515_o_0));
 INVx1_ASAP7_75t_R n_8516 (.A(n_8512_o_0),
    .Y(n_8516_o_0));
 AOI21xp33_ASAP7_75t_R n_8517 (.A1(n_8406_o_0),
    .A2(n_8478_o_0),
    .B(n_8381_o_0),
    .Y(n_8517_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8518 (.A1(n_8516_o_0),
    .A2(n_8510_o_0),
    .B(n_8517_o_0),
    .C(n_8426_o_0),
    .Y(n_8518_o_0));
 NAND3xp33_ASAP7_75t_R n_8519 (.A(n_8405_o_0),
    .B(n_8304_o_0),
    .C(n_8365_o_0),
    .Y(n_8519_o_0));
 NAND2xp33_ASAP7_75t_R n_852 (.A(n_849_o_0),
    .B(n_851_o_0),
    .Y(n_852_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8520 (.A1(n_8357_o_0),
    .A2(n_8400_o_0),
    .B(n_8519_o_0),
    .C(n_8427_o_0),
    .Y(n_8520_o_0));
 NAND2xp33_ASAP7_75t_R n_8521 (.A(n_8357_o_0),
    .B(n_8434_o_0),
    .Y(n_8521_o_0));
 AOI31xp33_ASAP7_75t_R n_8522 (.A1(n_8332_o_0),
    .A2(n_8345_o_0),
    .A3(n_8318_o_0),
    .B(n_8357_o_0),
    .Y(n_8522_o_0));
 OAI211xp5_ASAP7_75t_R n_8523 (.A1(n_8384_o_0),
    .A2(n_8370_o_0),
    .B(n_8385_o_0),
    .C(n_8365_o_0),
    .Y(n_8523_o_0));
 AOI21xp33_ASAP7_75t_R n_8524 (.A1(n_8522_o_0),
    .A2(n_8523_o_0),
    .B(n_8380_o_0),
    .Y(n_8524_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8525 (.A1(n_8521_o_0),
    .A2(net73),
    .B(n_8524_o_0),
    .C(n_8413_o_0),
    .Y(n_8525_o_0));
 OAI211xp5_ASAP7_75t_R n_8526 (.A1(n_8393_o_0),
    .A2(n_8520_o_0),
    .B(n_8525_o_0),
    .C(n_8441_o_0),
    .Y(n_8526_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8527 (.A1(n_8380_o_0),
    .A2(n_8508_o_0),
    .B(n_8518_o_0),
    .C(n_8526_o_0),
    .Y(n_8527_o_0));
 AOI211xp5_ASAP7_75t_R n_8528 (.A1(n_8505_o_0),
    .A2(n_8446_o_0),
    .B(n_8515_o_0),
    .C(n_8527_o_0),
    .Y(n_8528_o_0));
 NAND2xp33_ASAP7_75t_R n_8529 (.A(net73),
    .B(net38),
    .Y(n_8529_o_0));
 INVx1_ASAP7_75t_R n_853 (.A(_00909_),
    .Y(n_853_o_0));
 INVx1_ASAP7_75t_R n_8530 (.A(n_8470_o_0),
    .Y(n_8530_o_0));
 OAI21xp33_ASAP7_75t_R n_8531 (.A1(n_8318_o_0),
    .A2(n_8405_o_0),
    .B(n_8304_o_0),
    .Y(n_8531_o_0));
 NOR2xp33_ASAP7_75t_R n_8532 (.A(n_8530_o_0),
    .B(n_8531_o_0),
    .Y(n_8532_o_0));
 AOI31xp33_ASAP7_75t_R n_8533 (.A1(n_8446_o_0),
    .A2(n_8358_o_0),
    .A3(n_8529_o_0),
    .B(n_8532_o_0),
    .Y(n_8533_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8534 (.A1(n_8345_o_0),
    .A2(n_8318_o_0),
    .B(n_8434_o_0),
    .C(n_8408_o_0),
    .Y(n_8534_o_0));
 INVx1_ASAP7_75t_R n_8535 (.A(n_8534_o_0),
    .Y(n_8535_o_0));
 OAI21xp33_ASAP7_75t_R n_8536 (.A1(n_8383_o_0),
    .A2(n_8416_o_0),
    .B(n_8442_o_0),
    .Y(n_8536_o_0));
 NAND2xp33_ASAP7_75t_R n_8537 (.A(n_8304_o_0),
    .B(n_8431_o_0),
    .Y(n_8537_o_0));
 AOI31xp33_ASAP7_75t_R n_8538 (.A1(n_8384_o_0),
    .A2(n_8345_o_0),
    .A3(n_8318_o_0),
    .B(n_8357_o_0),
    .Y(n_8538_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8539 (.A1(n_8405_o_0),
    .A2(net73),
    .B(n_8538_o_0),
    .C(n_8446_o_0),
    .Y(n_8539_o_0));
 NAND2xp33_ASAP7_75t_R n_854 (.A(n_853_o_0),
    .B(n_850_o_0),
    .Y(n_854_o_0));
 OAI21xp33_ASAP7_75t_R n_8540 (.A1(n_8537_o_0),
    .A2(n_8349_o_0),
    .B(n_8539_o_0),
    .Y(n_8540_o_0));
 OAI211xp5_ASAP7_75t_R n_8541 (.A1(n_8535_o_0),
    .A2(n_8536_o_0),
    .B(n_8540_o_0),
    .C(n_8461_o_0),
    .Y(n_8541_o_0));
 OAI21xp33_ASAP7_75t_R n_8542 (.A1(n_8461_o_0),
    .A2(n_8533_o_0),
    .B(n_8541_o_0),
    .Y(n_8542_o_0));
 AOI21xp33_ASAP7_75t_R n_8543 (.A1(net67),
    .A2(n_8318_o_0),
    .B(n_8408_o_0),
    .Y(n_8543_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8544 (.A1(n_8365_o_0),
    .A2(n_8386_o_0),
    .B(n_8358_o_0),
    .C(n_8543_o_0),
    .Y(n_8544_o_0));
 INVx1_ASAP7_75t_R n_8545 (.A(n_8466_o_0),
    .Y(n_8545_o_0));
 NOR3xp33_ASAP7_75t_R n_8546 (.A(n_8346_o_0),
    .B(net73),
    .C(n_8357_o_0),
    .Y(n_8546_o_0));
 NOR5xp2_ASAP7_75t_R n_8547 (.A(n_8544_o_0),
    .B(n_8442_o_0),
    .C(n_8545_o_0),
    .D(n_8381_o_0),
    .E(n_8546_o_0),
    .Y(n_8547_o_0));
 OAI21xp33_ASAP7_75t_R n_8548 (.A1(n_8365_o_0),
    .A2(n_8346_o_0),
    .B(n_8304_o_0),
    .Y(n_8548_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8549 (.A1(_00905_),
    .A2(n_8287_o_0),
    .B(n_8288_o_0),
    .C(n_8380_o_0),
    .Y(n_8549_o_0));
 OAI21xp33_ASAP7_75t_R n_855 (.A1(n_850_o_0),
    .A2(n_853_o_0),
    .B(n_854_o_0),
    .Y(n_855_o_0));
 AOI21xp33_ASAP7_75t_R n_8550 (.A1(n_8522_o_0),
    .A2(n_8523_o_0),
    .B(n_8549_o_0),
    .Y(n_8550_o_0));
 OA21x2_ASAP7_75t_R n_8551 (.A1(n_8398_o_0),
    .A2(n_8548_o_0),
    .B(n_8550_o_0),
    .Y(n_8551_o_0));
 NAND5xp2_ASAP7_75t_R n_8552 (.A(n_8289_o_0),
    .B(n_8304_o_0),
    .C(n_8384_o_0),
    .D(net38),
    .E(net73),
    .Y(n_8552_o_0));
 NAND2xp33_ASAP7_75t_R n_8553 (.A(n_8318_o_0),
    .B(n_8370_o_0),
    .Y(n_8553_o_0));
 INVx1_ASAP7_75t_R n_8554 (.A(n_8553_o_0),
    .Y(n_8554_o_0));
 OAI211xp5_ASAP7_75t_R n_8555 (.A1(n_8435_o_0),
    .A2(n_8554_o_0),
    .B(n_8289_o_0),
    .C(n_8416_o_0),
    .Y(n_8555_o_0));
 INVx1_ASAP7_75t_R n_8556 (.A(n_8405_o_0),
    .Y(n_8556_o_0));
 OAI21xp33_ASAP7_75t_R n_8557 (.A1(net67),
    .A2(n_8365_o_0),
    .B(n_8357_o_0),
    .Y(n_8557_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8558 (.A1(n_8385_o_0),
    .A2(n_8389_o_0),
    .B(net73),
    .C(n_8408_o_0),
    .D(n_8289_o_0),
    .Y(n_8558_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8559 (.A1(n_8556_o_0),
    .A2(n_8365_o_0),
    .B(n_8557_o_0),
    .C(n_8558_o_0),
    .Y(n_8559_o_0));
 NAND2xp33_ASAP7_75t_R n_856 (.A(n_848_o_0),
    .B(n_855_o_0),
    .Y(n_856_o_0));
 AOI31xp33_ASAP7_75t_R n_8560 (.A1(n_8552_o_0),
    .A2(n_8555_o_0),
    .A3(n_8559_o_0),
    .B(n_8461_o_0),
    .Y(n_8560_o_0));
 NOR4xp25_ASAP7_75t_R n_8561 (.A(n_8547_o_0),
    .B(n_8551_o_0),
    .C(n_8560_o_0),
    .D(n_8295_o_0),
    .Y(n_8561_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8562 (.A1(n_8413_o_0),
    .A2(n_8542_o_0),
    .B(n_8561_o_0),
    .C(n_8279_o_0),
    .Y(n_8562_o_0));
 OAI21xp33_ASAP7_75t_R n_8563 (.A1(n_8279_o_0),
    .A2(n_8528_o_0),
    .B(n_8562_o_0),
    .Y(n_8563_o_0));
 AOI311xp33_ASAP7_75t_R n_8564 (.A1(n_8365_o_0),
    .A2(n_8389_o_0),
    .A3(n_8385_o_0),
    .B(n_8408_o_0),
    .C(n_8554_o_0),
    .Y(n_8564_o_0));
 AOI31xp33_ASAP7_75t_R n_8565 (.A1(n_8348_o_0),
    .A2(n_8358_o_0),
    .A3(n_8419_o_0),
    .B(n_8564_o_0),
    .Y(n_8565_o_0));
 AOI21xp33_ASAP7_75t_R n_8566 (.A1(net73),
    .A2(n_8434_o_0),
    .B(n_8408_o_0),
    .Y(n_8566_o_0));
 AOI21xp33_ASAP7_75t_R n_8567 (.A1(n_8492_o_0),
    .A2(n_8522_o_0),
    .B(n_8566_o_0),
    .Y(n_8567_o_0));
 OAI21xp33_ASAP7_75t_R n_8568 (.A1(n_8461_o_0),
    .A2(n_8567_o_0),
    .B(n_8295_o_0),
    .Y(n_8568_o_0));
 AOI21xp33_ASAP7_75t_R n_8569 (.A1(n_8385_o_0),
    .A2(n_8389_o_0),
    .B(n_8318_o_0),
    .Y(n_8569_o_0));
 NAND2xp33_ASAP7_75t_R n_857 (.A(key[17]),
    .B(ld),
    .Y(n_857_o_0));
 NOR2xp33_ASAP7_75t_R n_8570 (.A(n_8357_o_0),
    .B(n_8569_o_0),
    .Y(n_8570_o_0));
 NOR3xp33_ASAP7_75t_R n_8571 (.A(n_8464_o_0),
    .B(n_8408_o_0),
    .C(n_8430_o_0),
    .Y(n_8571_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8572 (.A1(n_8365_o_0),
    .A2(n_8386_o_0),
    .B(n_8570_o_0),
    .C(n_8571_o_0),
    .Y(n_8572_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8573 (.A1(net38),
    .A2(net73),
    .B(n_8384_o_0),
    .C(n_8304_o_0),
    .Y(n_8573_o_0));
 NAND3xp33_ASAP7_75t_R n_8574 (.A(n_8476_o_0),
    .B(n_8553_o_0),
    .C(n_8358_o_0),
    .Y(n_8574_o_0));
 AOI31xp33_ASAP7_75t_R n_8575 (.A1(n_8573_o_0),
    .A2(n_8574_o_0),
    .A3(n_8461_o_0),
    .B(n_8413_o_0),
    .Y(n_8575_o_0));
 OAI21xp33_ASAP7_75t_R n_8576 (.A1(n_8380_o_0),
    .A2(n_8572_o_0),
    .B(n_8575_o_0),
    .Y(n_8576_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8577 (.A1(n_8461_o_0),
    .A2(n_8565_o_0),
    .B(n_8568_o_0),
    .C(n_8576_o_0),
    .Y(n_8577_o_0));
 AOI211xp5_ASAP7_75t_R n_8578 (.A1(n_8399_o_0),
    .A2(n_8365_o_0),
    .B(n_8428_o_0),
    .C(n_8357_o_0),
    .Y(n_8578_o_0));
 AOI211xp5_ASAP7_75t_R n_8579 (.A1(n_8456_o_0),
    .A2(n_8474_o_0),
    .B(n_8578_o_0),
    .C(n_8380_o_0),
    .Y(n_8579_o_0));
 INVx1_ASAP7_75t_R n_858 (.A(n_857_o_0),
    .Y(n_858_o_0));
 AOI21xp33_ASAP7_75t_R n_8580 (.A1(n_8332_o_0),
    .A2(n_8345_o_0),
    .B(n_8365_o_0),
    .Y(n_8580_o_0));
 NAND2xp33_ASAP7_75t_R n_8581 (.A(n_8538_o_0),
    .B(n_8474_o_0),
    .Y(n_8581_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8582 (.A1(n_8510_o_0),
    .A2(n_8580_o_0),
    .B(n_8581_o_0),
    .C(n_8393_o_0),
    .Y(n_8582_o_0));
 NOR2xp33_ASAP7_75t_R n_8583 (.A(_00904_),
    .B(n_8379_o_0),
    .Y(n_8583_o_0));
 NOR2xp33_ASAP7_75t_R n_8584 (.A(n_8365_o_0),
    .B(n_8405_o_0),
    .Y(n_8584_o_0));
 OAI21xp33_ASAP7_75t_R n_8585 (.A1(n_8365_o_0),
    .A2(n_8399_o_0),
    .B(n_8419_o_0),
    .Y(n_8585_o_0));
 OAI32xp33_ASAP7_75t_R n_8586 (.A1(n_8408_o_0),
    .A2(n_8477_o_0),
    .A3(n_8584_o_0),
    .B1(n_8585_o_0),
    .B2(n_8357_o_0),
    .Y(n_8586_o_0));
 INVx1_ASAP7_75t_R n_8587 (.A(n_8392_o_0),
    .Y(n_8587_o_0));
 NAND3xp33_ASAP7_75t_R n_8588 (.A(n_8365_o_0),
    .B(net66),
    .C(n_8332_o_0),
    .Y(n_8588_o_0));
 OAI21xp33_ASAP7_75t_R n_8589 (.A1(n_8384_o_0),
    .A2(n_8365_o_0),
    .B(n_8345_o_0),
    .Y(n_8589_o_0));
 AOI31xp67_ASAP7_75t_R n_859 (.A1(n_827_o_0),
    .A2(n_852_o_0),
    .A3(n_856_o_0),
    .B(n_858_o_0),
    .Y(n_859_o_0));
 OAI22xp33_ASAP7_75t_R n_8590 (.A1(n_8588_o_0),
    .A2(n_8408_o_0),
    .B1(n_8589_o_0),
    .B2(n_8357_o_0),
    .Y(n_8590_o_0));
 AOI31xp33_ASAP7_75t_R n_8591 (.A1(net73),
    .A2(n_8357_o_0),
    .A3(n_8434_o_0),
    .B(n_8590_o_0),
    .Y(n_8591_o_0));
 OAI321xp33_ASAP7_75t_R n_8592 (.A1(n_8583_o_0),
    .A2(n_8586_o_0),
    .A3(n_8587_o_0),
    .B1(n_8461_o_0),
    .B2(n_8591_o_0),
    .C(n_8426_o_0),
    .Y(n_8592_o_0));
 OAI31xp33_ASAP7_75t_R n_8593 (.A1(n_8426_o_0),
    .A2(n_8579_o_0),
    .A3(n_8582_o_0),
    .B(n_8592_o_0),
    .Y(n_8593_o_0));
 OA22x2_ASAP7_75t_R n_8594 (.A1(n_8577_o_0),
    .A2(n_8446_o_0),
    .B1(n_8593_o_0),
    .B2(n_8441_o_0),
    .Y(n_8594_o_0));
 INVx1_ASAP7_75t_R n_8595 (.A(n_8347_o_0),
    .Y(n_8595_o_0));
 INVx1_ASAP7_75t_R n_8596 (.A(n_8450_o_0),
    .Y(n_8596_o_0));
 AOI21xp33_ASAP7_75t_R n_8597 (.A1(n_8570_o_0),
    .A2(n_8596_o_0),
    .B(n_8471_o_0),
    .Y(n_8597_o_0));
 AOI21xp33_ASAP7_75t_R n_8598 (.A1(n_8365_o_0),
    .A2(n_8332_o_0),
    .B(n_8357_o_0),
    .Y(n_8598_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8599 (.A1(n_8365_o_0),
    .A2(n_8405_o_0),
    .B(n_8598_o_0),
    .C(n_8393_o_0),
    .Y(n_8599_o_0));
 AND2x2_ASAP7_75t_R n_860 (.A(n_847_o_0),
    .B(n_859_o_0),
    .Y(n_860_o_0));
 OAI21xp33_ASAP7_75t_R n_8600 (.A1(n_8530_o_0),
    .A2(n_8531_o_0),
    .B(n_8599_o_0),
    .Y(n_8600_o_0));
 AOI21xp33_ASAP7_75t_R n_8601 (.A1(n_8295_o_0),
    .A2(n_8600_o_0),
    .B(n_8446_o_0),
    .Y(n_8601_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8602 (.A1(n_8595_o_0),
    .A2(n_8408_o_0),
    .B(n_8597_o_0),
    .C(n_8601_o_0),
    .Y(n_8602_o_0));
 NAND3xp33_ASAP7_75t_R n_8603 (.A(n_8431_o_0),
    .B(n_8553_o_0),
    .C(n_8358_o_0),
    .Y(n_8603_o_0));
 OAI31xp33_ASAP7_75t_R n_8604 (.A1(n_8357_o_0),
    .A2(n_8463_o_0),
    .A3(n_8390_o_0),
    .B(n_8381_o_0),
    .Y(n_8604_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8605 (.A1(n_8304_o_0),
    .A2(n_8453_o_0),
    .B(n_8604_o_0),
    .C(n_8414_o_0),
    .Y(n_8605_o_0));
 AOI31xp33_ASAP7_75t_R n_8606 (.A1(n_8603_o_0),
    .A2(n_8461_o_0),
    .A3(n_8475_o_0),
    .B(n_8605_o_0),
    .Y(n_8606_o_0));
 OAI21xp33_ASAP7_75t_R n_8607 (.A1(n_8602_o_0),
    .A2(n_8606_o_0),
    .B(n_8280_o_0),
    .Y(n_8607_o_0));
 INVx1_ASAP7_75t_R n_8608 (.A(n_8529_o_0),
    .Y(n_8608_o_0));
 NAND3xp33_ASAP7_75t_R n_8609 (.A(n_8474_o_0),
    .B(n_8418_o_0),
    .C(n_8358_o_0),
    .Y(n_8609_o_0));
 NOR2xp33_ASAP7_75t_R n_861 (.A(n_836_o_0),
    .B(n_860_o_0),
    .Y(n_861_o_0));
 OAI211xp5_ASAP7_75t_R n_8610 (.A1(n_8358_o_0),
    .A2(n_8608_o_0),
    .B(n_8609_o_0),
    .C(n_8393_o_0),
    .Y(n_8610_o_0));
 INVx1_ASAP7_75t_R n_8611 (.A(n_8485_o_0),
    .Y(n_8611_o_0));
 OAI21xp33_ASAP7_75t_R n_8612 (.A1(n_8365_o_0),
    .A2(n_8386_o_0),
    .B(n_8358_o_0),
    .Y(n_8612_o_0));
 AO21x1_ASAP7_75t_R n_8613 (.A1(n_8365_o_0),
    .A2(n_8371_o_0),
    .B(n_8612_o_0),
    .Y(n_8613_o_0));
 OAI31xp33_ASAP7_75t_R n_8614 (.A1(n_8408_o_0),
    .A2(n_8473_o_0),
    .A3(n_8611_o_0),
    .B(n_8613_o_0),
    .Y(n_8614_o_0));
 AOI21xp33_ASAP7_75t_R n_8615 (.A1(n_8380_o_0),
    .A2(n_8614_o_0),
    .B(n_8295_o_0),
    .Y(n_8615_o_0));
 AOI21xp33_ASAP7_75t_R n_8616 (.A1(n_8358_o_0),
    .A2(n_8454_o_0),
    .B(n_8566_o_0),
    .Y(n_8616_o_0));
 OAI31xp33_ASAP7_75t_R n_8617 (.A1(net38),
    .A2(n_8358_o_0),
    .A3(n_8365_o_0),
    .B(n_8380_o_0),
    .Y(n_8617_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8618 (.A1(n_8474_o_0),
    .A2(n_8538_o_0),
    .B(n_8617_o_0),
    .C(n_8413_o_0),
    .Y(n_8618_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8619 (.A1(n_8616_o_0),
    .A2(n_8393_o_0),
    .B(n_8618_o_0),
    .C(n_8446_o_0),
    .Y(n_8619_o_0));
 NOR2xp33_ASAP7_75t_R n_862 (.A(n_849_o_0),
    .B(n_851_o_0),
    .Y(n_862_o_0));
 AOI21xp33_ASAP7_75t_R n_8620 (.A1(n_8610_o_0),
    .A2(n_8615_o_0),
    .B(n_8619_o_0),
    .Y(n_8620_o_0));
 OAI22xp33_ASAP7_75t_R n_8621 (.A1(n_8594_o_0),
    .A2(n_8280_o_0),
    .B1(n_8607_o_0),
    .B2(n_8620_o_0),
    .Y(n_8621_o_0));
 NOR2xp33_ASAP7_75t_R n_8622 (.A(n_8506_o_0),
    .B(n_8455_o_0),
    .Y(n_8622_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8623 (.A1(n_8304_o_0),
    .A2(n_8470_o_0),
    .B(n_8622_o_0),
    .C(n_8474_o_0),
    .Y(n_8623_o_0));
 OAI21xp33_ASAP7_75t_R n_8624 (.A1(n_8358_o_0),
    .A2(n_8366_o_0),
    .B(n_8380_o_0),
    .Y(n_8624_o_0));
 INVx1_ASAP7_75t_R n_8625 (.A(n_8460_o_0),
    .Y(n_8625_o_0));
 AOI21xp33_ASAP7_75t_R n_8626 (.A1(n_8549_o_0),
    .A2(n_8624_o_0),
    .B(n_8625_o_0),
    .Y(n_8626_o_0));
 OAI21xp33_ASAP7_75t_R n_8627 (.A1(net66),
    .A2(n_8384_o_0),
    .B(n_8318_o_0),
    .Y(n_8627_o_0));
 AOI21xp33_ASAP7_75t_R n_8628 (.A1(n_8598_o_0),
    .A2(n_8627_o_0),
    .B(n_8441_o_0),
    .Y(n_8628_o_0));
 OAI21xp33_ASAP7_75t_R n_8629 (.A1(n_8569_o_0),
    .A2(n_8436_o_0),
    .B(n_8628_o_0),
    .Y(n_8629_o_0));
 NOR2xp33_ASAP7_75t_R n_863 (.A(n_848_o_0),
    .B(n_855_o_0),
    .Y(n_863_o_0));
 INVx1_ASAP7_75t_R n_8630 (.A(n_8464_o_0),
    .Y(n_8630_o_0));
 AOI31xp33_ASAP7_75t_R n_8631 (.A1(n_8304_o_0),
    .A2(n_8431_o_0),
    .A3(n_8630_o_0),
    .B(n_8446_o_0),
    .Y(n_8631_o_0));
 OAI21xp33_ASAP7_75t_R n_8632 (.A1(n_8588_o_0),
    .A2(n_8357_o_0),
    .B(n_8631_o_0),
    .Y(n_8632_o_0));
 AOI21xp33_ASAP7_75t_R n_8633 (.A1(n_8629_o_0),
    .A2(n_8632_o_0),
    .B(n_8380_o_0),
    .Y(n_8633_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8634 (.A1(n_8289_o_0),
    .A2(n_8623_o_0),
    .B(n_8626_o_0),
    .C(n_8633_o_0),
    .Y(n_8634_o_0));
 NAND2xp33_ASAP7_75t_R n_8635 (.A(n_8279_o_0),
    .B(n_8634_o_0),
    .Y(n_8635_o_0));
 INVx1_ASAP7_75t_R n_8636 (.A(n_8471_o_0),
    .Y(n_8636_o_0));
 AOI31xp33_ASAP7_75t_R n_8637 (.A1(n_8358_o_0),
    .A2(n_8492_o_0),
    .A3(n_8596_o_0),
    .B(n_8564_o_0),
    .Y(n_8637_o_0));
 NOR3xp33_ASAP7_75t_R n_8638 (.A(n_8569_o_0),
    .B(n_8554_o_0),
    .C(n_8357_o_0),
    .Y(n_8638_o_0));
 NOR2xp33_ASAP7_75t_R n_8639 (.A(n_8461_o_0),
    .B(n_8289_o_0),
    .Y(n_8639_o_0));
 OAI31xp33_ASAP7_75t_R n_864 (.A1(ld),
    .A2(n_862_o_0),
    .A3(n_863_o_0),
    .B(n_857_o_0),
    .Y(n_864_o_0));
 INVx1_ASAP7_75t_R n_8640 (.A(n_8639_o_0),
    .Y(n_8640_o_0));
 AOI21xp33_ASAP7_75t_R n_8641 (.A1(n_8447_o_0),
    .A2(n_8418_o_0),
    .B(n_8358_o_0),
    .Y(n_8641_o_0));
 OAI31xp33_ASAP7_75t_R n_8642 (.A1(n_8638_o_0),
    .A2(n_8640_o_0),
    .A3(n_8641_o_0),
    .B(n_8280_o_0),
    .Y(n_8642_o_0));
 AOI21xp33_ASAP7_75t_R n_8643 (.A1(n_8636_o_0),
    .A2(n_8637_o_0),
    .B(n_8642_o_0),
    .Y(n_8643_o_0));
 INVx1_ASAP7_75t_R n_8644 (.A(n_8536_o_0),
    .Y(n_8644_o_0));
 NOR2xp33_ASAP7_75t_R n_8645 (.A(n_8365_o_0),
    .B(n_8304_o_0),
    .Y(n_8645_o_0));
 NAND2xp33_ASAP7_75t_R n_8646 (.A(n_8386_o_0),
    .B(n_8645_o_0),
    .Y(n_8646_o_0));
 NOR2xp33_ASAP7_75t_R n_8647 (.A(net73),
    .B(n_8346_o_0),
    .Y(n_8647_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8648 (.A1(net67),
    .A2(net38),
    .B(net73),
    .C(n_8543_o_0),
    .Y(n_8648_o_0));
 OAI31xp33_ASAP7_75t_R n_8649 (.A1(n_8357_o_0),
    .A2(n_8390_o_0),
    .A3(n_8647_o_0),
    .B(n_8648_o_0),
    .Y(n_8649_o_0));
 OAI21xp33_ASAP7_75t_R n_865 (.A1(n_847_o_0),
    .A2(n_864_o_0),
    .B(n_836_o_0),
    .Y(n_865_o_0));
 OAI21xp33_ASAP7_75t_R n_8650 (.A1(n_8446_o_0),
    .A2(n_8649_o_0),
    .B(n_8380_o_0),
    .Y(n_8650_o_0));
 AO21x1_ASAP7_75t_R n_8651 (.A1(n_8644_o_0),
    .A2(n_8646_o_0),
    .B(n_8650_o_0),
    .Y(n_8651_o_0));
 AOI21xp33_ASAP7_75t_R n_8652 (.A1(n_8643_o_0),
    .A2(n_8651_o_0),
    .B(n_8414_o_0),
    .Y(n_8652_o_0));
 AOI21xp33_ASAP7_75t_R n_8653 (.A1(net67),
    .A2(net66),
    .B(n_8365_o_0),
    .Y(n_8653_o_0));
 INVx1_ASAP7_75t_R n_8654 (.A(n_8420_o_0),
    .Y(n_8654_o_0));
 OAI211xp5_ASAP7_75t_R n_8655 (.A1(n_8422_o_0),
    .A2(n_8653_o_0),
    .B(n_8654_o_0),
    .C(n_8380_o_0),
    .Y(n_8655_o_0));
 NOR2xp33_ASAP7_75t_R n_8656 (.A(net73),
    .B(n_8405_o_0),
    .Y(n_8656_o_0));
 AO21x1_ASAP7_75t_R n_8657 (.A1(net73),
    .A2(n_8434_o_0),
    .B(n_8423_o_0),
    .Y(n_8657_o_0));
 OAI31xp33_ASAP7_75t_R n_8658 (.A1(n_8408_o_0),
    .A2(n_8390_o_0),
    .A3(n_8656_o_0),
    .B(n_8657_o_0),
    .Y(n_8658_o_0));
 AOI21xp33_ASAP7_75t_R n_8659 (.A1(n_8393_o_0),
    .A2(n_8658_o_0),
    .B(n_8446_o_0),
    .Y(n_8659_o_0));
 INVx1_ASAP7_75t_R n_866 (.A(n_865_o_0),
    .Y(n_866_o_0));
 OAI211xp5_ASAP7_75t_R n_8660 (.A1(n_8386_o_0),
    .A2(net73),
    .B(n_8630_o_0),
    .C(n_8304_o_0),
    .Y(n_8660_o_0));
 OAI31xp33_ASAP7_75t_R n_8661 (.A1(n_8357_o_0),
    .A2(n_8400_o_0),
    .A3(n_8427_o_0),
    .B(n_8660_o_0),
    .Y(n_8661_o_0));
 OAI32xp33_ASAP7_75t_R n_8662 (.A1(n_8538_o_0),
    .A2(n_8641_o_0),
    .A3(n_8640_o_0),
    .B1(n_8661_o_0),
    .B2(n_8549_o_0),
    .Y(n_8662_o_0));
 AOI21xp33_ASAP7_75t_R n_8663 (.A1(n_8655_o_0),
    .A2(n_8659_o_0),
    .B(n_8662_o_0),
    .Y(n_8663_o_0));
 AOI211xp5_ASAP7_75t_R n_8664 (.A1(n_8630_o_0),
    .A2(n_8598_o_0),
    .B(n_8289_o_0),
    .C(n_8461_o_0),
    .Y(n_8664_o_0));
 OAI21xp33_ASAP7_75t_R n_8665 (.A1(n_8530_o_0),
    .A2(n_8531_o_0),
    .B(n_8664_o_0),
    .Y(n_8665_o_0));
 OAI311xp33_ASAP7_75t_R n_8666 (.A1(n_8289_o_0),
    .A2(n_8381_o_0),
    .A3(n_8573_o_0),
    .B1(n_8279_o_0),
    .C1(n_8665_o_0),
    .Y(n_8666_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8667 (.A1(net45),
    .A2(n_8365_o_0),
    .B(net67),
    .C(n_8358_o_0),
    .Y(n_8667_o_0));
 NAND3xp33_ASAP7_75t_R n_8668 (.A(n_8507_o_0),
    .B(n_8667_o_0),
    .C(n_8381_o_0),
    .Y(n_8668_o_0));
 AOI21xp33_ASAP7_75t_R n_8669 (.A1(n_8396_o_0),
    .A2(n_8476_o_0),
    .B(n_8304_o_0),
    .Y(n_8669_o_0));
 XOR2xp5_ASAP7_75t_R n_867 (.A(_00441_),
    .B(_00879_),
    .Y(n_867_o_0));
 INVx1_ASAP7_75t_R n_8670 (.A(n_8669_o_0),
    .Y(n_8670_o_0));
 OAI211xp5_ASAP7_75t_R n_8671 (.A1(n_8422_o_0),
    .A2(n_8580_o_0),
    .B(n_8670_o_0),
    .C(n_8380_o_0),
    .Y(n_8671_o_0));
 AOI21xp33_ASAP7_75t_R n_8672 (.A1(n_8668_o_0),
    .A2(n_8671_o_0),
    .B(n_8446_o_0),
    .Y(n_8672_o_0));
 OAI21xp33_ASAP7_75t_R n_8673 (.A1(n_8666_o_0),
    .A2(n_8672_o_0),
    .B(n_8426_o_0),
    .Y(n_8673_o_0));
 AOI21xp33_ASAP7_75t_R n_8674 (.A1(n_8280_o_0),
    .A2(n_8663_o_0),
    .B(n_8673_o_0),
    .Y(n_8674_o_0));
 AOI21xp33_ASAP7_75t_R n_8675 (.A1(n_8635_o_0),
    .A2(n_8652_o_0),
    .B(n_8674_o_0),
    .Y(n_8675_o_0));
 OAI31xp33_ASAP7_75t_R n_8676 (.A1(n_8365_o_0),
    .A2(n_8304_o_0),
    .A3(net38),
    .B(n_8393_o_0),
    .Y(n_8676_o_0));
 NOR3xp33_ASAP7_75t_R n_8677 (.A(n_8452_o_0),
    .B(n_8546_o_0),
    .C(n_8676_o_0),
    .Y(n_8677_o_0));
 AOI21xp33_ASAP7_75t_R n_8678 (.A1(n_8365_o_0),
    .A2(n_8434_o_0),
    .B(n_8304_o_0),
    .Y(n_8678_o_0));
 NAND2xp33_ASAP7_75t_R n_8679 (.A(net73),
    .B(net38),
    .Y(n_8679_o_0));
 INVx1_ASAP7_75t_R n_868 (.A(_00911_),
    .Y(n_868_o_0));
 OAI21xp33_ASAP7_75t_R n_8680 (.A1(n_8580_o_0),
    .A2(n_8510_o_0),
    .B(n_8380_o_0),
    .Y(n_8680_o_0));
 AOI21xp33_ASAP7_75t_R n_8681 (.A1(n_8678_o_0),
    .A2(n_8679_o_0),
    .B(n_8680_o_0),
    .Y(n_8681_o_0));
 NOR3xp33_ASAP7_75t_R n_8682 (.A(n_8677_o_0),
    .B(n_8681_o_0),
    .C(n_8441_o_0),
    .Y(n_8682_o_0));
 AOI211xp5_ASAP7_75t_R n_8683 (.A1(n_8455_o_0),
    .A2(n_8645_o_0),
    .B(n_8481_o_0),
    .C(n_8477_o_0),
    .Y(n_8683_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8684 (.A1(net45),
    .A2(net67),
    .B(net73),
    .C(n_8357_o_0),
    .Y(n_8684_o_0));
 INVx1_ASAP7_75t_R n_8685 (.A(n_8684_o_0),
    .Y(n_8685_o_0));
 AOI21xp33_ASAP7_75t_R n_8686 (.A1(n_8685_o_0),
    .A2(n_8391_o_0),
    .B(n_8465_o_0),
    .Y(n_8686_o_0));
 AOI211xp5_ASAP7_75t_R n_8687 (.A1(n_8380_o_0),
    .A2(n_8683_o_0),
    .B(n_8686_o_0),
    .C(n_8446_o_0),
    .Y(n_8687_o_0));
 AOI21xp33_ASAP7_75t_R n_8688 (.A1(n_8501_o_0),
    .A2(n_8401_o_0),
    .B(n_8358_o_0),
    .Y(n_8688_o_0));
 AOI31xp33_ASAP7_75t_R n_8689 (.A1(n_8358_o_0),
    .A2(n_8419_o_0),
    .A3(n_8630_o_0),
    .B(n_8688_o_0),
    .Y(n_8689_o_0));
 NAND2xp33_ASAP7_75t_R n_869 (.A(n_868_o_0),
    .B(n_867_o_0),
    .Y(n_869_o_0));
 OAI211xp5_ASAP7_75t_R n_8690 (.A1(n_8408_o_0),
    .A2(n_8556_o_0),
    .B(n_8612_o_0),
    .C(n_8381_o_0),
    .Y(n_8690_o_0));
 NAND2xp33_ASAP7_75t_R n_8691 (.A(n_8393_o_0),
    .B(n_8446_o_0),
    .Y(n_8691_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8692 (.A1(n_8466_o_0),
    .A2(n_8485_o_0),
    .B(n_8358_o_0),
    .C(n_8654_o_0),
    .D(n_8691_o_0),
    .Y(n_8692_o_0));
 NOR3xp33_ASAP7_75t_R n_8693 (.A(n_8464_o_0),
    .B(n_8400_o_0),
    .C(n_8357_o_0),
    .Y(n_8693_o_0));
 INVx1_ASAP7_75t_R n_8694 (.A(n_8693_o_0),
    .Y(n_8694_o_0));
 NAND3xp33_ASAP7_75t_R n_8695 (.A(n_8694_o_0),
    .B(n_8459_o_0),
    .C(n_8461_o_0),
    .Y(n_8695_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8696 (.A1(n_8441_o_0),
    .A2(n_8690_o_0),
    .B(n_8692_o_0),
    .C(n_8695_o_0),
    .Y(n_8696_o_0));
 OAI311xp33_ASAP7_75t_R n_8697 (.A1(n_8289_o_0),
    .A2(n_8381_o_0),
    .A3(n_8689_o_0),
    .B1(n_8279_o_0),
    .C1(n_8696_o_0),
    .Y(n_8697_o_0));
 OAI31xp33_ASAP7_75t_R n_8698 (.A1(n_8279_o_0),
    .A2(n_8682_o_0),
    .A3(n_8687_o_0),
    .B(n_8697_o_0),
    .Y(n_8698_o_0));
 INVx1_ASAP7_75t_R n_8699 (.A(n_8548_o_0),
    .Y(n_8699_o_0));
 OAI21xp33_ASAP7_75t_R n_870 (.A1(n_867_o_0),
    .A2(n_868_o_0),
    .B(n_869_o_0),
    .Y(n_870_o_0));
 OAI21xp33_ASAP7_75t_R n_8700 (.A1(n_8522_o_0),
    .A2(n_8699_o_0),
    .B(n_8380_o_0),
    .Y(n_8700_o_0));
 OAI21xp33_ASAP7_75t_R n_8701 (.A1(n_8365_o_0),
    .A2(n_8386_o_0),
    .B(n_8511_o_0),
    .Y(n_8701_o_0));
 AO21x1_ASAP7_75t_R n_8702 (.A1(n_8701_o_0),
    .A2(n_8409_o_0),
    .B(n_8380_o_0),
    .Y(n_8702_o_0));
 OAI21xp33_ASAP7_75t_R n_8703 (.A1(n_8358_o_0),
    .A2(n_8553_o_0),
    .B(n_8534_o_0),
    .Y(n_8703_o_0));
 OA21x2_ASAP7_75t_R n_8704 (.A1(n_8416_o_0),
    .A2(n_8427_o_0),
    .B(n_8442_o_0),
    .Y(n_8704_o_0));
 INVx1_ASAP7_75t_R n_8705 (.A(n_8549_o_0),
    .Y(n_8705_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8706 (.A1(n_8365_o_0),
    .A2(n_8357_o_0),
    .B(n_8704_o_0),
    .C(n_8705_o_0),
    .Y(n_8706_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8707 (.A1(n_8304_o_0),
    .A2(n_8347_o_0),
    .B(n_8703_o_0),
    .C(n_8461_o_0),
    .D(n_8706_o_0),
    .Y(n_8707_o_0));
 AOI31xp33_ASAP7_75t_R n_8708 (.A1(n_8441_o_0),
    .A2(n_8700_o_0),
    .A3(n_8702_o_0),
    .B(n_8707_o_0),
    .Y(n_8708_o_0));
 OAI22xp33_ASAP7_75t_R n_8709 (.A1(n_8484_o_0),
    .A2(net73),
    .B1(n_8464_o_0),
    .B2(n_8357_o_0),
    .Y(n_8709_o_0));
 NOR2xp33_ASAP7_75t_R n_871 (.A(_00943_),
    .B(n_870_o_0),
    .Y(n_871_o_0));
 OAI211xp5_ASAP7_75t_R n_8710 (.A1(net38),
    .A2(n_8365_o_0),
    .B(n_8431_o_0),
    .C(n_8358_o_0),
    .Y(n_8710_o_0));
 OAI211xp5_ASAP7_75t_R n_8711 (.A1(n_8349_o_0),
    .A2(n_8537_o_0),
    .B(n_8710_o_0),
    .C(n_8636_o_0),
    .Y(n_8711_o_0));
 OAI31xp33_ASAP7_75t_R n_8712 (.A1(n_8446_o_0),
    .A2(n_8393_o_0),
    .A3(n_8709_o_0),
    .B(n_8711_o_0),
    .Y(n_8712_o_0));
 INVx1_ASAP7_75t_R n_8713 (.A(n_8609_o_0),
    .Y(n_8713_o_0));
 AOI211xp5_ASAP7_75t_R n_8714 (.A1(net67),
    .A2(net73),
    .B(n_8357_o_0),
    .C(net45),
    .Y(n_8714_o_0));
 NOR2xp33_ASAP7_75t_R n_8715 (.A(n_8381_o_0),
    .B(n_8289_o_0),
    .Y(n_8715_o_0));
 OAI21xp33_ASAP7_75t_R n_8716 (.A1(n_8714_o_0),
    .A2(n_8688_o_0),
    .B(n_8715_o_0),
    .Y(n_8716_o_0));
 OAI31xp33_ASAP7_75t_R n_8717 (.A1(n_8461_o_0),
    .A2(n_8713_o_0),
    .A3(n_8536_o_0),
    .B(n_8716_o_0),
    .Y(n_8717_o_0));
 OAI31xp33_ASAP7_75t_R n_8718 (.A1(n_8279_o_0),
    .A2(n_8712_o_0),
    .A3(n_8717_o_0),
    .B(n_8414_o_0),
    .Y(n_8718_o_0));
 AOI21xp33_ASAP7_75t_R n_8719 (.A1(n_8279_o_0),
    .A2(n_8708_o_0),
    .B(n_8718_o_0),
    .Y(n_8719_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_872 (.A1(n_870_o_0),
    .A2(_00943_),
    .B(n_871_o_0),
    .C(_00975_),
    .Y(n_872_o_0));
 AOI21xp33_ASAP7_75t_R n_8720 (.A1(n_8295_o_0),
    .A2(n_8698_o_0),
    .B(n_8719_o_0),
    .Y(n_8720_o_0));
 NOR2xp33_ASAP7_75t_R n_8721 (.A(n_8473_o_0),
    .B(n_8548_o_0),
    .Y(n_8721_o_0));
 OAI21xp33_ASAP7_75t_R n_8722 (.A1(n_8408_o_0),
    .A2(n_8584_o_0),
    .B(n_8381_o_0),
    .Y(n_8722_o_0));
 AOI21xp33_ASAP7_75t_R n_8723 (.A1(n_8570_o_0),
    .A2(n_8485_o_0),
    .B(n_8722_o_0),
    .Y(n_8723_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8724 (.A1(n_8455_o_0),
    .A2(n_8645_o_0),
    .B(n_8721_o_0),
    .C(n_8461_o_0),
    .D(n_8723_o_0),
    .Y(n_8724_o_0));
 INVx1_ASAP7_75t_R n_8725 (.A(n_8688_o_0),
    .Y(n_8725_o_0));
 AOI21xp33_ASAP7_75t_R n_8726 (.A1(net38),
    .A2(n_8358_o_0),
    .B(n_8380_o_0),
    .Y(n_8726_o_0));
 INVx1_ASAP7_75t_R n_8727 (.A(n_8436_o_0),
    .Y(n_8727_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8728 (.A1(net67),
    .A2(net45),
    .B(net73),
    .C(n_8408_o_0),
    .Y(n_8728_o_0));
 OAI21xp33_ASAP7_75t_R n_8729 (.A1(n_8653_o_0),
    .A2(n_8728_o_0),
    .B(n_8380_o_0),
    .Y(n_8729_o_0));
 NAND2xp33_ASAP7_75t_R n_873 (.A(_00943_),
    .B(n_870_o_0),
    .Y(n_873_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8730 (.A1(n_8727_o_0),
    .A2(n_8501_o_0),
    .B(n_8729_o_0),
    .C(n_8441_o_0),
    .Y(n_8730_o_0));
 AOI21xp33_ASAP7_75t_R n_8731 (.A1(n_8725_o_0),
    .A2(n_8726_o_0),
    .B(n_8730_o_0),
    .Y(n_8731_o_0));
 AOI211xp5_ASAP7_75t_R n_8732 (.A1(n_8724_o_0),
    .A2(n_8446_o_0),
    .B(n_8731_o_0),
    .C(n_8414_o_0),
    .Y(n_8732_o_0));
 AOI21xp33_ASAP7_75t_R n_8733 (.A1(n_8422_o_0),
    .A2(n_8670_o_0),
    .B(n_8380_o_0),
    .Y(n_8733_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8734 (.A1(n_8450_o_0),
    .A2(n_8511_o_0),
    .B(n_8461_o_0),
    .C(n_8733_o_0),
    .Y(n_8734_o_0));
 OAI211xp5_ASAP7_75t_R n_8735 (.A1(n_8399_o_0),
    .A2(net73),
    .B(n_8630_o_0),
    .C(n_8304_o_0),
    .Y(n_8735_o_0));
 OAI31xp33_ASAP7_75t_R n_8736 (.A1(net67),
    .A2(n_8357_o_0),
    .A3(n_8450_o_0),
    .B(n_8735_o_0),
    .Y(n_8736_o_0));
 INVx1_ASAP7_75t_R n_8737 (.A(n_8580_o_0),
    .Y(n_8737_o_0));
 INVx1_ASAP7_75t_R n_8738 (.A(n_8404_o_0),
    .Y(n_8738_o_0));
 AOI21xp33_ASAP7_75t_R n_8739 (.A1(n_8737_o_0),
    .A2(n_8487_o_0),
    .B(n_8738_o_0),
    .Y(n_8739_o_0));
 INVx1_ASAP7_75t_R n_874 (.A(_00975_),
    .Y(n_874_o_0));
 NAND3xp33_ASAP7_75t_R n_8740 (.A(n_8739_o_0),
    .B(n_8441_o_0),
    .C(n_8381_o_0),
    .Y(n_8740_o_0));
 OAI31xp33_ASAP7_75t_R n_8741 (.A1(n_8381_o_0),
    .A2(n_8442_o_0),
    .A3(n_8736_o_0),
    .B(n_8740_o_0),
    .Y(n_8741_o_0));
 AOI211xp5_ASAP7_75t_R n_8742 (.A1(n_8734_o_0),
    .A2(n_8446_o_0),
    .B(n_8295_o_0),
    .C(n_8741_o_0),
    .Y(n_8742_o_0));
 INVx1_ASAP7_75t_R n_8743 (.A(n_8598_o_0),
    .Y(n_8743_o_0));
 OAI21xp33_ASAP7_75t_R n_8744 (.A1(n_8428_o_0),
    .A2(n_8531_o_0),
    .B(n_8743_o_0),
    .Y(n_8744_o_0));
 OAI211xp5_ASAP7_75t_R n_8745 (.A1(n_8304_o_0),
    .A2(n_8580_o_0),
    .B(n_8480_o_0),
    .C(n_8380_o_0),
    .Y(n_8745_o_0));
 OAI21xp33_ASAP7_75t_R n_8746 (.A1(n_8461_o_0),
    .A2(n_8744_o_0),
    .B(n_8745_o_0),
    .Y(n_8746_o_0));
 AOI211xp5_ASAP7_75t_R n_8747 (.A1(_00900_),
    .A2(n_8327_o_0),
    .B(net66),
    .C(n_8331_o_0),
    .Y(n_8747_o_0));
 OAI311xp33_ASAP7_75t_R n_8748 (.A1(net73),
    .A2(n_8747_o_0),
    .A3(n_8364_o_0),
    .B1(n_8627_o_0),
    .C1(n_8304_o_0),
    .Y(n_8748_o_0));
 OAI31xp33_ASAP7_75t_R n_8749 (.A1(n_8357_o_0),
    .A2(n_8569_o_0),
    .A3(n_8530_o_0),
    .B(n_8748_o_0),
    .Y(n_8749_o_0));
 OAI211xp5_ASAP7_75t_R n_875 (.A1(n_870_o_0),
    .A2(_00943_),
    .B(n_873_o_0),
    .C(n_874_o_0),
    .Y(n_875_o_0));
 AOI21xp33_ASAP7_75t_R n_8750 (.A1(n_8371_o_0),
    .A2(n_8358_o_0),
    .B(n_8441_o_0),
    .Y(n_8750_o_0));
 AOI22xp33_ASAP7_75t_R n_8751 (.A1(n_8446_o_0),
    .A2(n_8380_o_0),
    .B1(n_8531_o_0),
    .B2(n_8750_o_0),
    .Y(n_8751_o_0));
 AOI21xp33_ASAP7_75t_R n_8752 (.A1(n_8380_o_0),
    .A2(n_8749_o_0),
    .B(n_8751_o_0),
    .Y(n_8752_o_0));
 AOI211xp5_ASAP7_75t_R n_8753 (.A1(n_8746_o_0),
    .A2(n_8441_o_0),
    .B(n_8280_o_0),
    .C(n_8752_o_0),
    .Y(n_8753_o_0));
 OR2x2_ASAP7_75t_R n_8754 (.A(_00905_),
    .B(n_8286_o_0),
    .Y(n_8754_o_0));
 AOI31xp33_ASAP7_75t_R n_8755 (.A1(n_8365_o_0),
    .A2(net45),
    .A3(net67),
    .B(n_8408_o_0),
    .Y(n_8755_o_0));
 AOI21xp33_ASAP7_75t_R n_8756 (.A1(n_8429_o_0),
    .A2(n_8755_o_0),
    .B(n_8598_o_0),
    .Y(n_8756_o_0));
 NAND2xp33_ASAP7_75t_R n_8757 (.A(n_8318_o_0),
    .B(n_8357_o_0),
    .Y(n_8757_o_0));
 OAI21xp33_ASAP7_75t_R n_8758 (.A1(n_8399_o_0),
    .A2(n_8757_o_0),
    .B(n_8380_o_0),
    .Y(n_8758_o_0));
 AOI21xp33_ASAP7_75t_R n_8759 (.A1(n_8408_o_0),
    .A2(n_8737_o_0),
    .B(n_8758_o_0),
    .Y(n_8759_o_0));
 AND2x2_ASAP7_75t_R n_876 (.A(key[19]),
    .B(ld),
    .Y(n_876_o_0));
 AOI21xp33_ASAP7_75t_R n_8760 (.A1(n_8393_o_0),
    .A2(n_8756_o_0),
    .B(n_8759_o_0),
    .Y(n_8760_o_0));
 AOI311xp33_ASAP7_75t_R n_8761 (.A1(n_8365_o_0),
    .A2(n_8389_o_0),
    .A3(n_8385_o_0),
    .B(n_8408_o_0),
    .C(n_8427_o_0),
    .Y(n_8761_o_0));
 AOI31xp33_ASAP7_75t_R n_8762 (.A1(n_8358_o_0),
    .A2(n_8366_o_0),
    .A3(n_8470_o_0),
    .B(n_8761_o_0),
    .Y(n_8762_o_0));
 NOR2xp33_ASAP7_75t_R n_8763 (.A(n_8549_o_0),
    .B(n_8531_o_0),
    .Y(n_8763_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8764 (.A1(n_8358_o_0),
    .A2(n_8371_o_0),
    .B(n_8441_o_0),
    .C(n_8549_o_0),
    .D(n_8755_o_0),
    .Y(n_8764_o_0));
 OAI22xp33_ASAP7_75t_R n_8765 (.A1(n_8762_o_0),
    .A2(n_8381_o_0),
    .B1(n_8763_o_0),
    .B2(n_8764_o_0),
    .Y(n_8765_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8766 (.A1(n_8754_o_0),
    .A2(n_8440_o_0),
    .B(n_8760_o_0),
    .C(n_8765_o_0),
    .D(n_8280_o_0),
    .Y(n_8766_o_0));
 AOI311xp33_ASAP7_75t_R n_8767 (.A1(n_8365_o_0),
    .A2(net45),
    .A3(net67),
    .B(n_8408_o_0),
    .C(n_8427_o_0),
    .Y(n_8767_o_0));
 AOI31xp33_ASAP7_75t_R n_8768 (.A1(n_8358_o_0),
    .A2(n_8371_o_0),
    .A3(net73),
    .B(n_8767_o_0),
    .Y(n_8768_o_0));
 OAI32xp33_ASAP7_75t_R n_8769 (.A1(n_8537_o_0),
    .A2(n_8450_o_0),
    .A3(n_8461_o_0),
    .B1(n_8768_o_0),
    .B2(n_8381_o_0),
    .Y(n_8769_o_0));
 AOI31xp67_ASAP7_75t_R n_877 (.A1(n_827_o_0),
    .A2(n_872_o_0),
    .A3(n_875_o_0),
    .B(n_876_o_0),
    .Y(n_877_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8770 (.A1(n_8358_o_0),
    .A2(net67),
    .B(n_8417_o_0),
    .C(n_8381_o_0),
    .Y(n_8770_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8771 (.A1(n_8389_o_0),
    .A2(n_8385_o_0),
    .B(net73),
    .C(n_8538_o_0),
    .Y(n_8771_o_0));
 OAI31xp33_ASAP7_75t_R n_8772 (.A1(n_8408_o_0),
    .A2(n_8400_o_0),
    .A3(n_8464_o_0),
    .B(n_8771_o_0),
    .Y(n_8772_o_0));
 AOI21xp33_ASAP7_75t_R n_8773 (.A1(n_8380_o_0),
    .A2(n_8772_o_0),
    .B(n_8446_o_0),
    .Y(n_8773_o_0));
 AOI21xp33_ASAP7_75t_R n_8774 (.A1(n_8770_o_0),
    .A2(n_8773_o_0),
    .B(n_8295_o_0),
    .Y(n_8774_o_0));
 OAI21xp33_ASAP7_75t_R n_8775 (.A1(n_8482_o_0),
    .A2(n_8769_o_0),
    .B(n_8774_o_0),
    .Y(n_8775_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8776 (.A1(n_8753_o_0),
    .A2(n_8414_o_0),
    .B(n_8766_o_0),
    .C(n_8775_o_0),
    .Y(n_8776_o_0));
 OA31x2_ASAP7_75t_R n_8777 (.A1(n_8279_o_0),
    .A2(n_8732_o_0),
    .A3(n_8742_o_0),
    .B1(n_8776_o_0),
    .Y(n_8777_o_0));
 AOI211xp5_ASAP7_75t_R n_8778 (.A1(n_8434_o_0),
    .A2(n_8365_o_0),
    .B(n_8516_o_0),
    .C(n_8304_o_0),
    .Y(n_8778_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8779 (.A1(net73),
    .A2(n_8384_o_0),
    .B(n_8456_o_0),
    .C(n_8778_o_0),
    .Y(n_8779_o_0));
 AO31x2_ASAP7_75t_R n_878 (.A1(n_872_o_0),
    .A2(n_875_o_0),
    .A3(n_827_o_0),
    .B(n_876_o_0),
    .Y(n_878_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8780 (.A1(n_8365_o_0),
    .A2(net67),
    .B(net38),
    .C(n_8358_o_0),
    .Y(n_8780_o_0));
 AND3x1_ASAP7_75t_R n_8781 (.A(n_8372_o_0),
    .B(n_8780_o_0),
    .C(n_8461_o_0),
    .Y(n_8781_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8782 (.A1(n_8779_o_0),
    .A2(n_8381_o_0),
    .B(n_8781_o_0),
    .C(n_8442_o_0),
    .Y(n_8782_o_0));
 INVx1_ASAP7_75t_R n_8783 (.A(n_8538_o_0),
    .Y(n_8783_o_0));
 OAI22xp33_ASAP7_75t_R n_8784 (.A1(n_8611_o_0),
    .A2(n_8387_o_0),
    .B1(n_8400_o_0),
    .B2(n_8783_o_0),
    .Y(n_8784_o_0));
 AOI21xp33_ASAP7_75t_R n_8785 (.A1(n_8381_o_0),
    .A2(n_8784_o_0),
    .B(n_8442_o_0),
    .Y(n_8785_o_0));
 OAI21xp33_ASAP7_75t_R n_8786 (.A1(n_8616_o_0),
    .A2(n_8624_o_0),
    .B(n_8785_o_0),
    .Y(n_8786_o_0));
 AOI21xp33_ASAP7_75t_R n_8787 (.A1(net38),
    .A2(n_8365_o_0),
    .B(n_8408_o_0),
    .Y(n_8787_o_0));
 NAND2xp33_ASAP7_75t_R n_8788 (.A(net73),
    .B(net45),
    .Y(n_8788_o_0));
 OAI21xp33_ASAP7_75t_R n_8789 (.A1(net45),
    .A2(net73),
    .B(n_8788_o_0),
    .Y(n_8789_o_0));
 OAI21xp33_ASAP7_75t_R n_879 (.A1(n_841_o_0),
    .A2(n_837_o_0),
    .B(n_842_o_0),
    .Y(n_879_o_0));
 AOI22xp33_ASAP7_75t_R n_8790 (.A1(n_8787_o_0),
    .A2(n_8630_o_0),
    .B1(n_8358_o_0),
    .B2(n_8789_o_0),
    .Y(n_8790_o_0));
 INVx1_ASAP7_75t_R n_8791 (.A(n_8584_o_0),
    .Y(n_8791_o_0));
 AOI21xp33_ASAP7_75t_R n_8792 (.A1(n_8791_o_0),
    .A2(n_8570_o_0),
    .B(n_8393_o_0),
    .Y(n_8792_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8793 (.A1(net67),
    .A2(net73),
    .B(n_8408_o_0),
    .C(n_8792_o_0),
    .D(n_8442_o_0),
    .Y(n_8793_o_0));
 INVx1_ASAP7_75t_R n_8794 (.A(n_8578_o_0),
    .Y(n_8794_o_0));
 AOI32xp33_ASAP7_75t_R n_8795 (.A1(n_8358_o_0),
    .A2(n_8630_o_0),
    .A3(n_8401_o_0),
    .B1(n_8304_o_0),
    .B2(n_8470_o_0),
    .Y(n_8795_o_0));
 AOI21xp33_ASAP7_75t_R n_8796 (.A1(n_8715_o_0),
    .A2(n_8795_o_0),
    .B(n_8280_o_0),
    .Y(n_8796_o_0));
 OAI21xp33_ASAP7_75t_R n_8797 (.A1(n_8691_o_0),
    .A2(n_8794_o_0),
    .B(n_8796_o_0),
    .Y(n_8797_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8798 (.A1(n_8380_o_0),
    .A2(n_8790_o_0),
    .B(n_8793_o_0),
    .C(n_8797_o_0),
    .Y(n_8798_o_0));
 AOI31xp33_ASAP7_75t_R n_8799 (.A1(n_8280_o_0),
    .A2(n_8782_o_0),
    .A3(n_8786_o_0),
    .B(n_8798_o_0),
    .Y(n_8799_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_880 (.A1(n_879_o_0),
    .A2(ld),
    .B(n_845_o_0),
    .C(n_859_o_0),
    .Y(n_880_o_0));
 AOI31xp33_ASAP7_75t_R n_8800 (.A1(net73),
    .A2(n_8358_o_0),
    .A3(n_8384_o_0),
    .B(n_8441_o_0),
    .Y(n_8800_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8801 (.A1(n_8455_o_0),
    .A2(net73),
    .B(n_8416_o_0),
    .C(n_8800_o_0),
    .Y(n_8801_o_0));
 AOI21xp33_ASAP7_75t_R n_8802 (.A1(n_8304_o_0),
    .A2(n_8347_o_0),
    .B(n_8446_o_0),
    .Y(n_8802_o_0));
 OAI21xp33_ASAP7_75t_R n_8803 (.A1(n_8484_o_0),
    .A2(n_8506_o_0),
    .B(n_8802_o_0),
    .Y(n_8803_o_0));
 AOI21xp33_ASAP7_75t_R n_8804 (.A1(n_8801_o_0),
    .A2(n_8803_o_0),
    .B(n_8393_o_0),
    .Y(n_8804_o_0));
 NOR2xp33_ASAP7_75t_R n_8805 (.A(n_8318_o_0),
    .B(n_8484_o_0),
    .Y(n_8805_o_0));
 NOR2xp33_ASAP7_75t_R n_8806 (.A(n_8398_o_0),
    .B(n_8464_o_0),
    .Y(n_8806_o_0));
 AOI22xp33_ASAP7_75t_R n_8807 (.A1(n_8805_o_0),
    .A2(n_8358_o_0),
    .B1(n_8304_o_0),
    .B2(n_8806_o_0),
    .Y(n_8807_o_0));
 OAI21xp33_ASAP7_75t_R n_8808 (.A1(n_8506_o_0),
    .A2(n_8556_o_0),
    .B(n_8807_o_0),
    .Y(n_8808_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8809 (.A1(net67),
    .A2(net45),
    .B(n_8400_o_0),
    .C(n_8408_o_0),
    .Y(n_8809_o_0));
 INVx2_ASAP7_75t_R n_881 (.A(n_836_o_0),
    .Y(n_881_o_0));
 NAND2xp33_ASAP7_75t_R n_8810 (.A(net38),
    .B(n_8357_o_0),
    .Y(n_8810_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8811 (.A1(n_8809_o_0),
    .A2(n_8810_o_0),
    .B(n_8446_o_0),
    .C(n_8381_o_0),
    .Y(n_8811_o_0));
 AOI21xp33_ASAP7_75t_R n_8812 (.A1(n_8446_o_0),
    .A2(n_8808_o_0),
    .B(n_8811_o_0),
    .Y(n_8812_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8813 (.A1(n_8588_o_0),
    .A2(n_8357_o_0),
    .B(n_8804_o_0),
    .C(n_8812_o_0),
    .Y(n_8813_o_0));
 OAI211xp5_ASAP7_75t_R n_8814 (.A1(n_8365_o_0),
    .A2(n_8434_o_0),
    .B(n_8787_o_0),
    .C(n_8357_o_0),
    .Y(n_8814_o_0));
 NAND3xp33_ASAP7_75t_R n_8815 (.A(n_8418_o_0),
    .B(n_8447_o_0),
    .C(n_8358_o_0),
    .Y(n_8815_o_0));
 AOI211xp5_ASAP7_75t_R n_8816 (.A1(n_8814_o_0),
    .A2(n_8815_o_0),
    .B(n_8461_o_0),
    .C(n_8442_o_0),
    .Y(n_8816_o_0));
 INVx1_ASAP7_75t_R n_8817 (.A(n_8523_o_0),
    .Y(n_8817_o_0));
 AOI211xp5_ASAP7_75t_R n_8818 (.A1(n_8357_o_0),
    .A2(n_8817_o_0),
    .B(n_8691_o_0),
    .C(n_8669_o_0),
    .Y(n_8818_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8819 (.A1(n_8318_o_0),
    .A2(net38),
    .B(net67),
    .C(n_8304_o_0),
    .Y(n_8819_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_882 (.A1(n_847_o_0),
    .A2(n_859_o_0),
    .B(n_880_o_0),
    .C(n_881_o_0),
    .Y(n_882_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8820 (.A1(net45),
    .A2(net73),
    .B(n_8357_o_0),
    .C(n_8819_o_0),
    .Y(n_8820_o_0));
 NAND2xp33_ASAP7_75t_R n_8821 (.A(n_8441_o_0),
    .B(n_8447_o_0),
    .Y(n_8821_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8822 (.A1(n_8384_o_0),
    .A2(net38),
    .B(n_8357_o_0),
    .C(n_8684_o_0),
    .D(n_8821_o_0),
    .Y(n_8822_o_0));
 AOI211xp5_ASAP7_75t_R n_8823 (.A1(n_8446_o_0),
    .A2(n_8820_o_0),
    .B(n_8822_o_0),
    .C(n_8393_o_0),
    .Y(n_8823_o_0));
 NOR5xp2_ASAP7_75t_R n_8824 (.A(n_8816_o_0),
    .B(n_8818_o_0),
    .C(n_8295_o_0),
    .D(n_8280_o_0),
    .E(n_8823_o_0),
    .Y(n_8824_o_0));
 AOI31xp33_ASAP7_75t_R n_8825 (.A1(n_8280_o_0),
    .A2(n_8426_o_0),
    .A3(n_8813_o_0),
    .B(n_8824_o_0),
    .Y(n_8825_o_0));
 OAI21xp33_ASAP7_75t_R n_8826 (.A1(n_8426_o_0),
    .A2(n_8799_o_0),
    .B(n_8825_o_0),
    .Y(n_8826_o_0));
 NOR2xp33_ASAP7_75t_R n_8827 (.A(n_8464_o_0),
    .B(n_8743_o_0),
    .Y(n_8827_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8828 (.A1(n_8304_o_0),
    .A2(n_8474_o_0),
    .B(n_8827_o_0),
    .C(n_8791_o_0),
    .Y(n_8828_o_0));
 NOR3xp33_ASAP7_75t_R n_8829 (.A(n_8556_o_0),
    .B(n_8365_o_0),
    .C(n_8408_o_0),
    .Y(n_8829_o_0));
 NAND2xp33_ASAP7_75t_R n_883 (.A(n_878_o_0),
    .B(n_882_o_0),
    .Y(n_883_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8830 (.A1(n_8358_o_0),
    .A2(n_8470_o_0),
    .B(n_8829_o_0),
    .C(n_8523_o_0),
    .Y(n_8830_o_0));
 AOI21xp33_ASAP7_75t_R n_8831 (.A1(n_8304_o_0),
    .A2(n_8347_o_0),
    .B(n_8380_o_0),
    .Y(n_8831_o_0));
 AOI22xp33_ASAP7_75t_R n_8832 (.A1(n_8828_o_0),
    .A2(n_8461_o_0),
    .B1(n_8830_o_0),
    .B2(n_8831_o_0),
    .Y(n_8832_o_0));
 AOI211xp5_ASAP7_75t_R n_8833 (.A1(n_8408_o_0),
    .A2(n_8554_o_0),
    .B(n_8449_o_0),
    .C(n_8647_o_0),
    .Y(n_8833_o_0));
 OA211x2_ASAP7_75t_R n_8834 (.A1(n_8358_o_0),
    .A2(n_8399_o_0),
    .B(n_8809_o_0),
    .C(n_8380_o_0),
    .Y(n_8834_o_0));
 OAI31xp33_ASAP7_75t_R n_8835 (.A1(n_8441_o_0),
    .A2(n_8833_o_0),
    .A3(n_8834_o_0),
    .B(n_8414_o_0),
    .Y(n_8835_o_0));
 AOI21xp33_ASAP7_75t_R n_8836 (.A1(n_8289_o_0),
    .A2(n_8832_o_0),
    .B(n_8835_o_0),
    .Y(n_8836_o_0));
 NOR3xp33_ASAP7_75t_R n_8837 (.A(n_8477_o_0),
    .B(n_8390_o_0),
    .C(n_8408_o_0),
    .Y(n_8837_o_0));
 AOI21xp33_ASAP7_75t_R n_8838 (.A1(n_8358_o_0),
    .A2(n_8529_o_0),
    .B(n_8837_o_0),
    .Y(n_8838_o_0));
 NOR2xp33_ASAP7_75t_R n_8839 (.A(n_8400_o_0),
    .B(n_8436_o_0),
    .Y(n_8839_o_0));
 AOI21xp33_ASAP7_75t_R n_884 (.A1(net32),
    .A2(n_860_o_0),
    .B(n_883_o_0),
    .Y(n_884_o_0));
 AOI31xp33_ASAP7_75t_R n_8840 (.A1(n_8358_o_0),
    .A2(n_8391_o_0),
    .A3(n_8523_o_0),
    .B(n_8839_o_0),
    .Y(n_8840_o_0));
 OAI31xp33_ASAP7_75t_R n_8841 (.A1(n_8289_o_0),
    .A2(n_8840_o_0),
    .A3(n_8381_o_0),
    .B(n_8413_o_0),
    .Y(n_8841_o_0));
 INVx1_ASAP7_75t_R n_8842 (.A(n_8703_o_0),
    .Y(n_8842_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8843 (.A1(n_8358_o_0),
    .A2(n_8405_o_0),
    .B(n_8449_o_0),
    .C(n_8289_o_0),
    .Y(n_8843_o_0));
 AOI31xp33_ASAP7_75t_R n_8844 (.A1(n_8842_o_0),
    .A2(n_8461_o_0),
    .A3(n_8459_o_0),
    .B(n_8843_o_0),
    .Y(n_8844_o_0));
 AOI211xp5_ASAP7_75t_R n_8845 (.A1(n_8639_o_0),
    .A2(n_8838_o_0),
    .B(n_8841_o_0),
    .C(n_8844_o_0),
    .Y(n_8845_o_0));
 OAI21xp33_ASAP7_75t_R n_8846 (.A1(n_8421_o_0),
    .A2(n_8495_o_0),
    .B(n_8609_o_0),
    .Y(n_8846_o_0));
 NOR2xp33_ASAP7_75t_R n_8847 (.A(n_8430_o_0),
    .B(n_8383_o_0),
    .Y(n_8847_o_0));
 OAI21xp33_ASAP7_75t_R n_8848 (.A1(net67),
    .A2(n_8408_o_0),
    .B(n_8461_o_0),
    .Y(n_8848_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8849 (.A1(n_8847_o_0),
    .A2(n_8358_o_0),
    .B(n_8848_o_0),
    .C(n_8441_o_0),
    .Y(n_8849_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_885 (.A1(n_861_o_0),
    .A2(n_866_o_0),
    .B(n_877_o_0),
    .C(n_884_o_0),
    .Y(n_885_o_0));
 AOI21xp33_ASAP7_75t_R n_8850 (.A1(n_8381_o_0),
    .A2(n_8846_o_0),
    .B(n_8849_o_0),
    .Y(n_8850_o_0));
 INVx1_ASAP7_75t_R n_8851 (.A(n_8387_o_0),
    .Y(n_8851_o_0));
 OAI21xp33_ASAP7_75t_R n_8852 (.A1(n_8357_o_0),
    .A2(n_8463_o_0),
    .B(n_8705_o_0),
    .Y(n_8852_o_0));
 AOI21xp33_ASAP7_75t_R n_8853 (.A1(n_8851_o_0),
    .A2(n_8791_o_0),
    .B(n_8852_o_0),
    .Y(n_8853_o_0));
 AOI21xp33_ASAP7_75t_R n_8854 (.A1(n_8422_o_0),
    .A2(n_8728_o_0),
    .B(n_8640_o_0),
    .Y(n_8854_o_0));
 NOR3xp33_ASAP7_75t_R n_8855 (.A(n_8850_o_0),
    .B(n_8853_o_0),
    .C(n_8854_o_0),
    .Y(n_8855_o_0));
 OAI22xp33_ASAP7_75t_R n_8856 (.A1(n_8493_o_0),
    .A2(n_8357_o_0),
    .B1(n_8436_o_0),
    .B2(n_8569_o_0),
    .Y(n_8856_o_0));
 INVx1_ASAP7_75t_R n_8857 (.A(n_8806_o_0),
    .Y(n_8857_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8858 (.A1(n_8408_o_0),
    .A2(n_8857_o_0),
    .B(n_8603_o_0),
    .C(n_8691_o_0),
    .Y(n_8858_o_0));
 AOI21xp33_ASAP7_75t_R n_8859 (.A1(n_8715_o_0),
    .A2(n_8856_o_0),
    .B(n_8858_o_0),
    .Y(n_8859_o_0));
 NAND2xp33_ASAP7_75t_R n_886 (.A(n_864_o_0),
    .B(n_836_o_0),
    .Y(n_886_o_0));
 AOI31xp33_ASAP7_75t_R n_8860 (.A1(n_8358_o_0),
    .A2(n_8484_o_0),
    .A3(n_8365_o_0),
    .B(n_8393_o_0),
    .Y(n_8860_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8861 (.A1(n_8506_o_0),
    .A2(n_8556_o_0),
    .B(n_8860_o_0),
    .C(n_8727_o_0),
    .Y(n_8861_o_0));
 AOI31xp33_ASAP7_75t_R n_8862 (.A1(n_8434_o_0),
    .A2(n_8860_o_0),
    .A3(n_8365_o_0),
    .B(n_8436_o_0),
    .Y(n_8862_o_0));
 OAI321xp33_ASAP7_75t_R n_8863 (.A1(n_8685_o_0),
    .A2(n_8693_o_0),
    .A3(n_8380_o_0),
    .B1(n_8861_o_0),
    .B2(n_8862_o_0),
    .C(n_8441_o_0),
    .Y(n_8863_o_0));
 AOI31xp33_ASAP7_75t_R n_8864 (.A1(n_8426_o_0),
    .A2(n_8859_o_0),
    .A3(n_8863_o_0),
    .B(n_8280_o_0),
    .Y(n_8864_o_0));
 OAI21xp33_ASAP7_75t_R n_8865 (.A1(n_8414_o_0),
    .A2(n_8855_o_0),
    .B(n_8864_o_0),
    .Y(n_8865_o_0));
 OAI31xp33_ASAP7_75t_R n_8866 (.A1(n_8836_o_0),
    .A2(n_8845_o_0),
    .A3(n_8279_o_0),
    .B(n_8865_o_0),
    .Y(n_8866_o_0));
 XOR2xp5_ASAP7_75t_R n_8867 (.A(_01105_),
    .B(_01106_),
    .Y(n_8867_o_0));
 XNOR2xp5_ASAP7_75t_R n_8868 (.A(_01066_),
    .B(n_8867_o_0),
    .Y(n_8868_o_0));
 NOR2xp33_ASAP7_75t_R n_8869 (.A(n_4227_o_0),
    .B(n_8868_o_0),
    .Y(n_8869_o_0));
 INVx1_ASAP7_75t_R n_887 (.A(n_886_o_0),
    .Y(n_887_o_0));
 NOR2xp33_ASAP7_75t_R n_8870 (.A(_00699_),
    .B(net),
    .Y(n_8870_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8871 (.A1(n_4227_o_0),
    .A2(n_8868_o_0),
    .B(n_8869_o_0),
    .C(net),
    .D(n_8870_o_0),
    .Y(n_8871_o_0));
 XNOR2xp5_ASAP7_75t_R n_8872 (.A(n_1342_o_0),
    .B(n_8871_o_0),
    .Y(n_8872_o_0));
 INVx1_ASAP7_75t_R n_8873 (.A(n_8872_o_0),
    .Y(n_8873_o_0));
 XNOR2xp5_ASAP7_75t_R n_8874 (.A(_01105_),
    .B(n_4298_o_0),
    .Y(n_8874_o_0));
 NOR2xp33_ASAP7_75t_R n_8875 (.A(n_4394_o_0),
    .B(n_8874_o_0),
    .Y(n_8875_o_0));
 NOR2xp33_ASAP7_75t_R n_8876 (.A(_00700_),
    .B(net),
    .Y(n_8876_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8877 (.A1(n_4394_o_0),
    .A2(n_8874_o_0),
    .B(n_8875_o_0),
    .C(net),
    .D(n_8876_o_0),
    .Y(n_8877_o_0));
 NOR2xp33_ASAP7_75t_R n_8878 (.A(_00938_),
    .B(n_8877_o_0),
    .Y(n_8878_o_0));
 AND2x2_ASAP7_75t_R n_8879 (.A(_00938_),
    .B(n_8877_o_0),
    .Y(n_8879_o_0));
 NAND2xp33_ASAP7_75t_R n_888 (.A(n_847_o_0),
    .B(n_859_o_0),
    .Y(n_888_o_0));
 NOR2xp33_ASAP7_75t_R n_8880 (.A(n_8878_o_0),
    .B(n_8879_o_0),
    .Y(n_8880_o_0));
 XOR2xp5_ASAP7_75t_R n_8881 (.A(_01102_),
    .B(_01106_),
    .Y(n_8881_o_0));
 XNOR2xp5_ASAP7_75t_R n_8882 (.A(n_4296_o_0),
    .B(n_8881_o_0),
    .Y(n_8882_o_0));
 XNOR2xp5_ASAP7_75t_R n_8883 (.A(_01103_),
    .B(n_6568_o_0),
    .Y(n_8883_o_0));
 NAND2xp33_ASAP7_75t_R n_8884 (.A(n_8883_o_0),
    .B(n_8882_o_0),
    .Y(n_8884_o_0));
 OAI21xp33_ASAP7_75t_R n_8885 (.A1(n_8882_o_0),
    .A2(n_8883_o_0),
    .B(n_8884_o_0),
    .Y(n_8885_o_0));
 NOR2xp33_ASAP7_75t_R n_8886 (.A(_00702_),
    .B(net77),
    .Y(n_8886_o_0));
 AOI21xp33_ASAP7_75t_R n_8887 (.A1(net),
    .A2(n_8885_o_0),
    .B(n_8886_o_0),
    .Y(n_8887_o_0));
 NAND2xp33_ASAP7_75t_R n_8888 (.A(_00936_),
    .B(n_8887_o_0),
    .Y(n_8888_o_0));
 OAI21xp33_ASAP7_75t_R n_8889 (.A1(_00936_),
    .A2(n_8887_o_0),
    .B(n_8888_o_0),
    .Y(n_8889_o_0));
 OAI21xp33_ASAP7_75t_R n_889 (.A1(n_847_o_0),
    .A2(n_859_o_0),
    .B(n_888_o_0),
    .Y(n_889_o_0));
 XOR2xp5_ASAP7_75t_R n_8890 (.A(_01099_),
    .B(_01106_),
    .Y(n_8890_o_0));
 NAND2xp33_ASAP7_75t_R n_8891 (.A(n_6574_o_0),
    .B(n_8890_o_0),
    .Y(n_8891_o_0));
 OAI21xp33_ASAP7_75t_R n_8892 (.A1(n_6574_o_0),
    .A2(n_8890_o_0),
    .B(n_8891_o_0),
    .Y(n_8892_o_0));
 NAND2xp33_ASAP7_75t_R n_8893 (.A(_01100_),
    .B(n_4185_o_0),
    .Y(n_8893_o_0));
 OAI21xp33_ASAP7_75t_R n_8894 (.A1(_01100_),
    .A2(n_4185_o_0),
    .B(n_8893_o_0),
    .Y(n_8894_o_0));
 NAND2xp33_ASAP7_75t_R n_8895 (.A(n_8894_o_0),
    .B(n_8892_o_0),
    .Y(n_8895_o_0));
 OAI211xp5_ASAP7_75t_R n_8896 (.A1(n_8892_o_0),
    .A2(n_8894_o_0),
    .B(n_8895_o_0),
    .C(net39),
    .Y(n_8896_o_0));
 NAND2xp33_ASAP7_75t_R n_8897 (.A(_00593_),
    .B(n_3021_o_0),
    .Y(n_8897_o_0));
 INVx1_ASAP7_75t_R n_8898 (.A(_00933_),
    .Y(n_8898_o_0));
 OAI21xp33_ASAP7_75t_R n_8899 (.A1(n_8894_o_0),
    .A2(n_8892_o_0),
    .B(net39),
    .Y(n_8899_o_0));
 OAI21xp33_ASAP7_75t_R n_890 (.A1(n_836_o_0),
    .A2(n_889_o_0),
    .B(n_877_o_0),
    .Y(n_890_o_0));
 XNOR2xp5_ASAP7_75t_R n_8900 (.A(_01099_),
    .B(_01106_),
    .Y(n_8900_o_0));
 XNOR2xp5_ASAP7_75t_R n_8901 (.A(n_8900_o_0),
    .B(n_6574_o_0),
    .Y(n_8901_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8902 (.A1(_01100_),
    .A2(n_4185_o_0),
    .B(n_8893_o_0),
    .C(n_8901_o_0),
    .Y(n_8902_o_0));
 OAI311xp33_ASAP7_75t_R n_8903 (.A1(n_3021_o_0),
    .A2(n_8899_o_0),
    .A3(n_8902_o_0),
    .B1(n_8898_o_0),
    .C1(n_8897_o_0),
    .Y(n_8903_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8904 (.A1(n_8896_o_0),
    .A2(n_8897_o_0),
    .B(n_8898_o_0),
    .C(n_8903_o_0),
    .Y(n_8904_o_0));
 XOR2xp5_ASAP7_75t_R n_8905 (.A(_01052_),
    .B(_01067_),
    .Y(n_8905_o_0));
 NAND2xp33_ASAP7_75t_R n_8906 (.A(_01012_),
    .B(n_8905_o_0),
    .Y(n_8906_o_0));
 OAI21xp33_ASAP7_75t_R n_8907 (.A1(_01012_),
    .A2(n_8905_o_0),
    .B(n_8906_o_0),
    .Y(n_8907_o_0));
 OAI211xp5_ASAP7_75t_R n_8908 (.A1(_01012_),
    .A2(n_8905_o_0),
    .B(n_8906_o_0),
    .C(n_8890_o_0),
    .Y(n_8908_o_0));
 INVx1_ASAP7_75t_R n_8909 (.A(n_8908_o_0),
    .Y(n_8909_o_0));
 INVx1_ASAP7_75t_R n_891 (.A(n_829_o_0),
    .Y(n_891_o_0));
 NOR2xp33_ASAP7_75t_R n_8910 (.A(_00594_),
    .B(net77),
    .Y(n_8910_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8911 (.A1(n_8900_o_0),
    .A2(n_8907_o_0),
    .B(n_8909_o_0),
    .C(net39),
    .D(n_8910_o_0),
    .Y(n_8911_o_0));
 NAND2xp33_ASAP7_75t_R n_8912 (.A(n_8900_o_0),
    .B(n_8907_o_0),
    .Y(n_8912_o_0));
 INVx1_ASAP7_75t_R n_8913 (.A(n_8910_o_0),
    .Y(n_8913_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8914 (.A1(n_8908_o_0),
    .A2(n_8912_o_0),
    .B(net3),
    .C(n_8913_o_0),
    .D(_00932_),
    .Y(n_8914_o_0));
 AOI21x1_ASAP7_75t_R n_8915 (.A1(_00932_),
    .A2(n_8911_o_0),
    .B(n_8914_o_0),
    .Y(n_8915_o_0));
 XOR2xp5_ASAP7_75t_R n_8916 (.A(_01014_),
    .B(_01054_),
    .Y(n_8916_o_0));
 INVx1_ASAP7_75t_R n_8917 (.A(_01101_),
    .Y(n_8917_o_0));
 NAND2xp33_ASAP7_75t_R n_8918 (.A(n_8917_o_0),
    .B(n_8916_o_0),
    .Y(n_8918_o_0));
 OAI21xp33_ASAP7_75t_R n_8919 (.A1(n_8916_o_0),
    .A2(n_8917_o_0),
    .B(n_8918_o_0),
    .Y(n_8919_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_892 (.A1(n_847_o_0),
    .A2(n_859_o_0),
    .B(n_888_o_0),
    .C(n_881_o_0),
    .Y(n_892_o_0));
 NOR2xp33_ASAP7_75t_R n_8920 (.A(n_8917_o_0),
    .B(n_8916_o_0),
    .Y(n_8920_o_0));
 AOI211xp5_ASAP7_75t_R n_8921 (.A1(n_8916_o_0),
    .A2(n_8917_o_0),
    .B(n_8920_o_0),
    .C(n_6589_o_0),
    .Y(n_8921_o_0));
 NOR2xp33_ASAP7_75t_R n_8922 (.A(_00596_),
    .B(_00858_),
    .Y(n_8922_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8923 (.A1(n_6589_o_0),
    .A2(n_8919_o_0),
    .B(n_8921_o_0),
    .C(net77),
    .D(n_8922_o_0),
    .Y(n_8923_o_0));
 INVx1_ASAP7_75t_R n_8924 (.A(_00934_),
    .Y(n_8924_o_0));
 NAND2xp33_ASAP7_75t_R n_8925 (.A(n_8924_o_0),
    .B(n_8923_o_0),
    .Y(n_8925_o_0));
 OAI21x1_ASAP7_75t_R n_8926 (.A1(n_8923_o_0),
    .A2(n_8924_o_0),
    .B(n_8925_o_0),
    .Y(n_8926_o_0));
 AOI21xp33_ASAP7_75t_R n_8927 (.A1(net48),
    .A2(n_8915_o_0),
    .B(n_8926_o_0),
    .Y(n_8927_o_0));
 INVx1_ASAP7_75t_R n_8928 (.A(n_8927_o_0),
    .Y(n_8928_o_0));
 XNOR2xp5_ASAP7_75t_R n_8929 (.A(_01102_),
    .B(n_6616_o_0),
    .Y(n_8929_o_0));
 NOR2xp33_ASAP7_75t_R n_893 (.A(n_877_o_0),
    .B(n_892_o_0),
    .Y(n_893_o_0));
 XNOR2xp5_ASAP7_75t_R n_8930 (.A(_01015_),
    .B(_01055_),
    .Y(n_8930_o_0));
 XNOR2xp5_ASAP7_75t_R n_8931 (.A(_01101_),
    .B(_01106_),
    .Y(n_8931_o_0));
 XNOR2xp5_ASAP7_75t_R n_8932 (.A(n_8930_o_0),
    .B(n_8931_o_0),
    .Y(n_8932_o_0));
 XOR2xp5_ASAP7_75t_R n_8933 (.A(n_8929_o_0),
    .B(n_8932_o_0),
    .Y(n_8933_o_0));
 NOR2xp33_ASAP7_75t_R n_8934 (.A(_00703_),
    .B(net77),
    .Y(n_8934_o_0));
 AOI21xp33_ASAP7_75t_R n_8935 (.A1(net77),
    .A2(n_8933_o_0),
    .B(n_8934_o_0),
    .Y(n_8935_o_0));
 XNOR2xp5_ASAP7_75t_R n_8936 (.A(n_8929_o_0),
    .B(n_8932_o_0),
    .Y(n_8936_o_0));
 OR2x2_ASAP7_75t_R n_8937 (.A(_00703_),
    .B(net77),
    .Y(n_8937_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8938 (.A1(net1),
    .A2(n_8936_o_0),
    .B(n_8937_o_0),
    .C(_00935_),
    .Y(n_8938_o_0));
 AOI21x1_ASAP7_75t_R n_8939 (.A1(_00935_),
    .A2(n_8935_o_0),
    .B(n_8938_o_0),
    .Y(n_8939_o_0));
 NOR2xp33_ASAP7_75t_R n_894 (.A(n_891_o_0),
    .B(n_893_o_0),
    .Y(n_894_o_0));
 OAI21xp33_ASAP7_75t_R n_8940 (.A1(net9),
    .A2(n_8936_o_0),
    .B(n_8937_o_0),
    .Y(n_8940_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8941 (.A1(n_8933_o_0),
    .A2(net),
    .B(n_8934_o_0),
    .C(_00935_),
    .Y(n_8941_o_0));
 OAI21xp5_ASAP7_75t_R n_8942 (.A1(_00935_),
    .A2(n_8940_o_0),
    .B(n_8941_o_0),
    .Y(n_8942_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8943 (.A1(n_8896_o_0),
    .A2(n_8897_o_0),
    .B(n_8898_o_0),
    .C(n_8903_o_0),
    .D(n_8915_o_0),
    .Y(n_8943_o_0));
 AOI211xp5_ASAP7_75t_R n_8944 (.A1(_00932_),
    .A2(n_8911_o_0),
    .B(n_8904_o_0),
    .C(n_8914_o_0),
    .Y(n_8944_o_0));
 OAI21xp33_ASAP7_75t_R n_8945 (.A1(n_8943_o_0),
    .A2(n_8944_o_0),
    .B(n_8926_o_0),
    .Y(n_8945_o_0));
 AO21x1_ASAP7_75t_R n_8946 (.A1(_00932_),
    .A2(n_8911_o_0),
    .B(n_8914_o_0),
    .Y(n_8946_o_0));
 XNOR2x1_ASAP7_75t_R n_8947 (.B(n_8923_o_0),
    .Y(n_8947_o_0),
    .A(_00934_));
 NAND3xp33_ASAP7_75t_R n_8948 (.A(n_8946_o_0),
    .B(net19),
    .C(n_8947_o_0),
    .Y(n_8948_o_0));
 AOI211xp5_ASAP7_75t_R n_8949 (.A1(n_8946_o_0),
    .A2(net48),
    .B(n_8939_o_0),
    .C(n_8947_o_0),
    .Y(n_8949_o_0));
 XOR2xp5_ASAP7_75t_R n_895 (.A(_00443_),
    .B(_00881_),
    .Y(n_895_o_0));
 AOI31xp33_ASAP7_75t_R n_8950 (.A1(n_8942_o_0),
    .A2(n_8945_o_0),
    .A3(n_8948_o_0),
    .B(n_8949_o_0),
    .Y(n_8950_o_0));
 OAI21xp33_ASAP7_75t_R n_8951 (.A1(n_8928_o_0),
    .A2(n_8939_o_0),
    .B(n_8950_o_0),
    .Y(n_8951_o_0));
 NOR2xp33_ASAP7_75t_R n_8952 (.A(n_8904_o_0),
    .B(n_8926_o_0),
    .Y(n_8952_o_0));
 INVx1_ASAP7_75t_R n_8953 (.A(n_8952_o_0),
    .Y(n_8953_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8954 (.A1(_00932_),
    .A2(n_8911_o_0),
    .B(n_8914_o_0),
    .C(n_8904_o_0),
    .Y(n_8954_o_0));
 INVx1_ASAP7_75t_R n_8955 (.A(n_8896_o_0),
    .Y(n_8955_o_0));
 INVx1_ASAP7_75t_R n_8956 (.A(n_8897_o_0),
    .Y(n_8956_o_0));
 AO21x1_ASAP7_75t_R n_8957 (.A1(n_8896_o_0),
    .A2(n_8897_o_0),
    .B(n_8898_o_0),
    .Y(n_8957_o_0));
 OAI311xp33_ASAP7_75t_R n_8958 (.A1(_00933_),
    .A2(n_8955_o_0),
    .A3(n_8956_o_0),
    .B1(n_8915_o_0),
    .C1(n_8957_o_0),
    .Y(n_8958_o_0));
 AOI31xp33_ASAP7_75t_R n_8959 (.A1(n_8954_o_0),
    .A2(n_8958_o_0),
    .A3(n_8926_o_0),
    .B(n_8939_o_0),
    .Y(n_8959_o_0));
 XOR2xp5_ASAP7_75t_R n_896 (.A(_00913_),
    .B(n_895_o_0),
    .Y(n_896_o_0));
 OAI21xp33_ASAP7_75t_R n_8960 (.A1(n_8946_o_0),
    .A2(n_8904_o_0),
    .B(n_8954_o_0),
    .Y(n_8960_o_0));
 INVx1_ASAP7_75t_R n_8961 (.A(_00935_),
    .Y(n_8961_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_8962 (.A1(n_8933_o_0),
    .A2(net),
    .B(n_8934_o_0),
    .C(n_8961_o_0),
    .Y(n_8962_o_0));
 OAI21xp5_ASAP7_75t_R n_8963 (.A1(n_8961_o_0),
    .A2(n_8940_o_0),
    .B(n_8962_o_0),
    .Y(n_8963_o_0));
 AOI21xp33_ASAP7_75t_R n_8964 (.A1(n_8947_o_0),
    .A2(n_8960_o_0),
    .B(n_8963_o_0),
    .Y(n_8964_o_0));
 AOI211xp5_ASAP7_75t_R n_8965 (.A1(n_8953_o_0),
    .A2(n_8959_o_0),
    .B(n_8964_o_0),
    .C(n_8889_o_0),
    .Y(n_8965_o_0));
 AOI21xp33_ASAP7_75t_R n_8966 (.A1(n_8889_o_0),
    .A2(n_8951_o_0),
    .B(n_8965_o_0),
    .Y(n_8966_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_8967 (.A1(net1),
    .A2(n_8936_o_0),
    .B(n_8937_o_0),
    .C(n_8961_o_0),
    .Y(n_8967_o_0));
 AOI21x1_ASAP7_75t_R n_8968 (.A1(n_8961_o_0),
    .A2(n_8935_o_0),
    .B(n_8967_o_0),
    .Y(n_8968_o_0));
 NOR3xp33_ASAP7_75t_R n_8969 (.A(n_8946_o_0),
    .B(net48),
    .C(n_8947_o_0),
    .Y(n_8969_o_0));
 NOR2xp33_ASAP7_75t_R n_897 (.A(_00945_),
    .B(n_896_o_0),
    .Y(n_897_o_0));
 NOR2xp33_ASAP7_75t_R n_8970 (.A(n_8926_o_0),
    .B(n_8915_o_0),
    .Y(n_8970_o_0));
 AOI211xp5_ASAP7_75t_R n_8971 (.A1(n_8885_o_0),
    .A2(net39),
    .B(_00936_),
    .C(n_8886_o_0),
    .Y(n_8971_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8972 (.A1(n_8885_o_0),
    .A2(net),
    .B(n_8886_o_0),
    .C(_00936_),
    .D(n_8971_o_0),
    .Y(n_8972_o_0));
 OAI31xp33_ASAP7_75t_R n_8973 (.A1(n_8968_o_0),
    .A2(n_8969_o_0),
    .A3(n_8970_o_0),
    .B(n_8972_o_0),
    .Y(n_8973_o_0));
 INVx1_ASAP7_75t_R n_8974 (.A(n_8904_o_0),
    .Y(n_8974_o_0));
 AOI211xp5_ASAP7_75t_R n_8975 (.A1(n_8915_o_0),
    .A2(n_8926_o_0),
    .B(n_8974_o_0),
    .C(n_8942_o_0),
    .Y(n_8975_o_0));
 NOR3xp33_ASAP7_75t_R n_8976 (.A(n_8915_o_0),
    .B(n_8926_o_0),
    .C(n_8904_o_0),
    .Y(n_8976_o_0));
 NAND2xp33_ASAP7_75t_R n_8977 (.A(net48),
    .B(n_8926_o_0),
    .Y(n_8977_o_0));
 INVx1_ASAP7_75t_R n_8978 (.A(n_8977_o_0),
    .Y(n_8978_o_0));
 OAI21xp33_ASAP7_75t_R n_8979 (.A1(net48),
    .A2(n_8946_o_0),
    .B(n_8926_o_0),
    .Y(n_8979_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_898 (.A1(n_896_o_0),
    .A2(_00945_),
    .B(n_897_o_0),
    .C(_00977_),
    .Y(n_898_o_0));
 NOR2xp33_ASAP7_75t_R n_8980 (.A(n_8968_o_0),
    .B(n_8970_o_0),
    .Y(n_8980_o_0));
 AOI21xp33_ASAP7_75t_R n_8981 (.A1(n_8979_o_0),
    .A2(n_8980_o_0),
    .B(n_8889_o_0),
    .Y(n_8981_o_0));
 OAI31xp33_ASAP7_75t_R n_8982 (.A1(n_8939_o_0),
    .A2(n_8976_o_0),
    .A3(n_8978_o_0),
    .B(n_8981_o_0),
    .Y(n_8982_o_0));
 XNOR2xp5_ASAP7_75t_R n_8983 (.A(_00938_),
    .B(n_8877_o_0),
    .Y(n_8983_o_0));
 INVx1_ASAP7_75t_R n_8984 (.A(n_8983_o_0),
    .Y(n_8984_o_0));
 OAI211xp5_ASAP7_75t_R n_8985 (.A1(n_8973_o_0),
    .A2(n_8975_o_0),
    .B(n_8982_o_0),
    .C(n_8984_o_0),
    .Y(n_8985_o_0));
 OAI21xp33_ASAP7_75t_R n_8986 (.A1(n_8880_o_0),
    .A2(n_8966_o_0),
    .B(n_8985_o_0),
    .Y(n_8986_o_0));
 NAND2xp33_ASAP7_75t_R n_8987 (.A(n_4266_o_0),
    .B(n_4338_o_0),
    .Y(n_8987_o_0));
 OAI21xp33_ASAP7_75t_R n_8988 (.A1(n_4266_o_0),
    .A2(n_4338_o_0),
    .B(n_8987_o_0),
    .Y(n_8988_o_0));
 NOR2xp33_ASAP7_75t_R n_8989 (.A(_01104_),
    .B(n_8988_o_0),
    .Y(n_8989_o_0));
 NAND2xp33_ASAP7_75t_R n_899 (.A(_00945_),
    .B(n_896_o_0),
    .Y(n_899_o_0));
 NOR2xp33_ASAP7_75t_R n_8990 (.A(_00701_),
    .B(net),
    .Y(n_8990_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_8991 (.A1(n_8988_o_0),
    .A2(_01104_),
    .B(n_8989_o_0),
    .C(net),
    .D(n_8990_o_0),
    .Y(n_8991_o_0));
 XNOR2xp5_ASAP7_75t_R n_8992 (.A(_00937_),
    .B(n_8991_o_0),
    .Y(n_8992_o_0));
 INVx1_ASAP7_75t_R n_8993 (.A(n_8992_o_0),
    .Y(n_8993_o_0));
 NAND2xp33_ASAP7_75t_R n_8994 (.A(n_8926_o_0),
    .B(n_8915_o_0),
    .Y(n_8994_o_0));
 NAND2xp33_ASAP7_75t_R n_8995 (.A(net48),
    .B(n_8946_o_0),
    .Y(n_8995_o_0));
 AOI21xp33_ASAP7_75t_R n_8996 (.A1(n_8994_o_0),
    .A2(n_8995_o_0),
    .B(n_8963_o_0),
    .Y(n_8996_o_0));
 NOR2xp33_ASAP7_75t_R n_8997 (.A(n_8972_o_0),
    .B(n_8996_o_0),
    .Y(n_8997_o_0));
 OAI21xp33_ASAP7_75t_R n_8998 (.A1(n_8947_o_0),
    .A2(n_8946_o_0),
    .B(n_8963_o_0),
    .Y(n_8998_o_0));
 INVx1_ASAP7_75t_R n_8999 (.A(n_8998_o_0),
    .Y(n_8999_o_0));
 INVx1_ASAP7_75t_R n_900 (.A(_00977_),
    .Y(n_900_o_0));
 NAND2xp33_ASAP7_75t_R n_9000 (.A(n_8995_o_0),
    .B(n_8999_o_0),
    .Y(n_9000_o_0));
 NAND3xp33_ASAP7_75t_R n_9001 (.A(n_8915_o_0),
    .B(n_8926_o_0),
    .C(n_8904_o_0),
    .Y(n_9001_o_0));
 NOR3xp33_ASAP7_75t_R n_9002 (.A(n_8974_o_0),
    .B(n_8926_o_0),
    .C(n_8915_o_0),
    .Y(n_9002_o_0));
 NOR2xp33_ASAP7_75t_R n_9003 (.A(n_8968_o_0),
    .B(n_9002_o_0),
    .Y(n_9003_o_0));
 NAND3xp33_ASAP7_75t_R n_9004 (.A(n_8974_o_0),
    .B(n_8947_o_0),
    .C(n_8915_o_0),
    .Y(n_9004_o_0));
 INVx1_ASAP7_75t_R n_9005 (.A(n_9004_o_0),
    .Y(n_9005_o_0));
 AOI21xp33_ASAP7_75t_R n_9006 (.A1(n_8954_o_0),
    .A2(n_8958_o_0),
    .B(n_8947_o_0),
    .Y(n_9006_o_0));
 OAI31xp33_ASAP7_75t_R n_9007 (.A1(n_8939_o_0),
    .A2(n_9005_o_0),
    .A3(n_9006_o_0),
    .B(n_8972_o_0),
    .Y(n_9007_o_0));
 INVx1_ASAP7_75t_R n_9008 (.A(n_8880_o_0),
    .Y(n_9008_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9009 (.A1(n_9001_o_0),
    .A2(n_9003_o_0),
    .B(n_9007_o_0),
    .C(n_9008_o_0),
    .Y(n_9009_o_0));
 OAI211xp5_ASAP7_75t_R n_901 (.A1(n_896_o_0),
    .A2(_00945_),
    .B(n_899_o_0),
    .C(n_900_o_0),
    .Y(n_901_o_0));
 INVx1_ASAP7_75t_R n_9010 (.A(n_8972_o_0),
    .Y(n_9010_o_0));
 OAI21xp33_ASAP7_75t_R n_9011 (.A1(n_8926_o_0),
    .A2(n_8915_o_0),
    .B(n_8968_o_0),
    .Y(n_9011_o_0));
 NOR2xp33_ASAP7_75t_R n_9012 (.A(n_8904_o_0),
    .B(n_8915_o_0),
    .Y(n_9012_o_0));
 OAI21xp33_ASAP7_75t_R n_9013 (.A1(n_8947_o_0),
    .A2(n_9012_o_0),
    .B(n_8939_o_0),
    .Y(n_9013_o_0));
 AOI21xp33_ASAP7_75t_R n_9014 (.A1(n_9011_o_0),
    .A2(n_9013_o_0),
    .B(n_8976_o_0),
    .Y(n_9014_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9015 (.A1(n_8958_o_0),
    .A2(n_8954_o_0),
    .B(n_8947_o_0),
    .C(n_8942_o_0),
    .Y(n_9015_o_0));
 AOI21xp33_ASAP7_75t_R n_9016 (.A1(n_8915_o_0),
    .A2(n_8974_o_0),
    .B(n_8926_o_0),
    .Y(n_9016_o_0));
 AOI21xp33_ASAP7_75t_R n_9017 (.A1(n_8946_o_0),
    .A2(n_8926_o_0),
    .B(n_8939_o_0),
    .Y(n_9017_o_0));
 NAND3xp33_ASAP7_75t_R n_9018 (.A(n_8974_o_0),
    .B(n_8946_o_0),
    .C(n_8947_o_0),
    .Y(n_9018_o_0));
 AOI21xp33_ASAP7_75t_R n_9019 (.A1(n_9017_o_0),
    .A2(n_9018_o_0),
    .B(n_8889_o_0),
    .Y(n_9019_o_0));
 AND2x2_ASAP7_75t_R n_902 (.A(key[21]),
    .B(ld),
    .Y(n_902_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9020 (.A1(n_9015_o_0),
    .A2(n_9016_o_0),
    .B(n_9019_o_0),
    .C(n_8983_o_0),
    .Y(n_9020_o_0));
 OAI21xp33_ASAP7_75t_R n_9021 (.A1(n_9010_o_0),
    .A2(n_9014_o_0),
    .B(n_9020_o_0),
    .Y(n_9021_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9022 (.A1(n_8997_o_0),
    .A2(n_9000_o_0),
    .B(n_9009_o_0),
    .C(n_9021_o_0),
    .Y(n_9022_o_0));
 NAND2xp33_ASAP7_75t_R n_9023 (.A(_00937_),
    .B(n_8991_o_0),
    .Y(n_9023_o_0));
 OAI21xp33_ASAP7_75t_R n_9024 (.A1(_00937_),
    .A2(n_8991_o_0),
    .B(n_9023_o_0),
    .Y(n_9024_o_0));
 OAI22xp33_ASAP7_75t_R n_9025 (.A1(n_8986_o_0),
    .A2(n_8993_o_0),
    .B1(n_9022_o_0),
    .B2(n_9024_o_0),
    .Y(n_9025_o_0));
 AOI21xp33_ASAP7_75t_R n_9026 (.A1(n_9001_o_0),
    .A2(n_9018_o_0),
    .B(n_8942_o_0),
    .Y(n_9026_o_0));
 AOI21xp33_ASAP7_75t_R n_9027 (.A1(n_8926_o_0),
    .A2(n_8960_o_0),
    .B(n_8963_o_0),
    .Y(n_9027_o_0));
 OAI31xp33_ASAP7_75t_R n_9028 (.A1(net64),
    .A2(n_9026_o_0),
    .A3(n_9027_o_0),
    .B(n_8880_o_0),
    .Y(n_9028_o_0));
 INVx1_ASAP7_75t_R n_9029 (.A(n_9012_o_0),
    .Y(n_9029_o_0));
 AOI31xp67_ASAP7_75t_R n_903 (.A1(n_827_o_0),
    .A2(n_898_o_0),
    .A3(n_901_o_0),
    .B(n_902_o_0),
    .Y(n_903_o_0));
 INVx1_ASAP7_75t_R n_9030 (.A(n_8973_o_0),
    .Y(n_9030_o_0));
 OAI31xp33_ASAP7_75t_R n_9031 (.A1(n_8926_o_0),
    .A2(n_9029_o_0),
    .A3(n_8939_o_0),
    .B(n_9030_o_0),
    .Y(n_9031_o_0));
 INVx1_ASAP7_75t_R n_9032 (.A(n_9031_o_0),
    .Y(n_9032_o_0));
 NAND2xp33_ASAP7_75t_R n_9033 (.A(n_8904_o_0),
    .B(n_8926_o_0),
    .Y(n_9033_o_0));
 INVx1_ASAP7_75t_R n_9034 (.A(n_9033_o_0),
    .Y(n_9034_o_0));
 AOI31xp33_ASAP7_75t_R n_9035 (.A1(n_8954_o_0),
    .A2(n_8958_o_0),
    .A3(n_8947_o_0),
    .B(n_8939_o_0),
    .Y(n_9035_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9036 (.A1(n_8947_o_0),
    .A2(n_9034_o_0),
    .B(n_8942_o_0),
    .C(n_9035_o_0),
    .Y(n_9036_o_0));
 OA21x2_ASAP7_75t_R n_9037 (.A1(_00936_),
    .A2(n_8887_o_0),
    .B(n_8888_o_0),
    .Y(n_9037_o_0));
 AOI21xp33_ASAP7_75t_R n_9038 (.A1(n_8968_o_0),
    .A2(n_9002_o_0),
    .B(n_9037_o_0),
    .Y(n_9038_o_0));
 AOI21xp33_ASAP7_75t_R n_9039 (.A1(net48),
    .A2(n_8946_o_0),
    .B(n_8947_o_0),
    .Y(n_9039_o_0));
 INVx1_ASAP7_75t_R n_904 (.A(n_903_o_0),
    .Y(n_904_o_0));
 NAND2xp33_ASAP7_75t_R n_9040 (.A(n_8915_o_0),
    .B(n_8947_o_0),
    .Y(n_9040_o_0));
 INVx1_ASAP7_75t_R n_9041 (.A(n_9040_o_0),
    .Y(n_9041_o_0));
 OAI21xp33_ASAP7_75t_R n_9042 (.A1(n_9039_o_0),
    .A2(n_9041_o_0),
    .B(n_8939_o_0),
    .Y(n_9042_o_0));
 NAND3xp33_ASAP7_75t_R n_9043 (.A(n_8974_o_0),
    .B(n_8926_o_0),
    .C(n_8946_o_0),
    .Y(n_9043_o_0));
 OAI211xp5_ASAP7_75t_R n_9044 (.A1(n_9012_o_0),
    .A2(n_8926_o_0),
    .B(n_9043_o_0),
    .C(n_8968_o_0),
    .Y(n_9044_o_0));
 AOI31xp33_ASAP7_75t_R n_9045 (.A1(n_9038_o_0),
    .A2(n_9042_o_0),
    .A3(n_9044_o_0),
    .B(n_8984_o_0),
    .Y(n_9045_o_0));
 INVx1_ASAP7_75t_R n_9046 (.A(n_9024_o_0),
    .Y(n_9046_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9047 (.A1(net64),
    .A2(n_9036_o_0),
    .B(n_9045_o_0),
    .C(n_9046_o_0),
    .Y(n_9047_o_0));
 OAI21xp33_ASAP7_75t_R n_9048 (.A1(n_9028_o_0),
    .A2(n_9032_o_0),
    .B(n_9047_o_0),
    .Y(n_9048_o_0));
 NOR3xp33_ASAP7_75t_R n_9049 (.A(n_8974_o_0),
    .B(n_8926_o_0),
    .C(n_8946_o_0),
    .Y(n_9049_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_905 (.A1(n_887_o_0),
    .A2(n_890_o_0),
    .B(n_894_o_0),
    .C(n_904_o_0),
    .Y(n_905_o_0));
 INVx1_ASAP7_75t_R n_9050 (.A(n_9049_o_0),
    .Y(n_9050_o_0));
 NAND2xp33_ASAP7_75t_R n_9051 (.A(net48),
    .B(n_8946_o_0),
    .Y(n_9051_o_0));
 OAI31xp33_ASAP7_75t_R n_9052 (.A1(n_8947_o_0),
    .A2(n_9051_o_0),
    .A3(n_8963_o_0),
    .B(n_9010_o_0),
    .Y(n_9052_o_0));
 AOI31xp33_ASAP7_75t_R n_9053 (.A1(n_8963_o_0),
    .A2(n_9050_o_0),
    .A3(n_9043_o_0),
    .B(n_9052_o_0),
    .Y(n_9053_o_0));
 NOR2xp33_ASAP7_75t_R n_9054 (.A(n_8915_o_0),
    .B(n_8974_o_0),
    .Y(n_9054_o_0));
 NOR2xp33_ASAP7_75t_R n_9055 (.A(n_8947_o_0),
    .B(n_8942_o_0),
    .Y(n_9055_o_0));
 NOR3xp33_ASAP7_75t_R n_9056 (.A(n_8947_o_0),
    .B(n_8915_o_0),
    .C(net19),
    .Y(n_9056_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9057 (.A1(n_8915_o_0),
    .A2(net19),
    .B(n_8926_o_0),
    .C(n_8939_o_0),
    .Y(n_9057_o_0));
 OAI21xp33_ASAP7_75t_R n_9058 (.A1(n_9056_o_0),
    .A2(n_9057_o_0),
    .B(n_8889_o_0),
    .Y(n_9058_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9059 (.A1(n_9054_o_0),
    .A2(n_9055_o_0),
    .B(n_9058_o_0),
    .C(n_8983_o_0),
    .Y(n_9059_o_0));
 OAI21xp33_ASAP7_75t_R n_906 (.A1(net16),
    .A2(n_885_o_0),
    .B(n_905_o_0),
    .Y(n_906_o_0));
 AOI21xp33_ASAP7_75t_R n_9060 (.A1(net48),
    .A2(n_8946_o_0),
    .B(n_8926_o_0),
    .Y(n_9060_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9061 (.A1(n_9054_o_0),
    .A2(n_8926_o_0),
    .B(n_9060_o_0),
    .C(n_8968_o_0),
    .Y(n_9061_o_0));
 NAND3xp33_ASAP7_75t_R n_9062 (.A(n_9061_o_0),
    .B(n_9013_o_0),
    .C(n_9010_o_0),
    .Y(n_9062_o_0));
 OAI21xp33_ASAP7_75t_R n_9063 (.A1(n_8915_o_0),
    .A2(n_8947_o_0),
    .B(n_8939_o_0),
    .Y(n_9063_o_0));
 OAI21xp33_ASAP7_75t_R n_9064 (.A1(n_8947_o_0),
    .A2(net19),
    .B(n_9035_o_0),
    .Y(n_9064_o_0));
 OAI211xp5_ASAP7_75t_R n_9065 (.A1(n_9063_o_0),
    .A2(n_9049_o_0),
    .B(n_9064_o_0),
    .C(n_8889_o_0),
    .Y(n_9065_o_0));
 AOI31xp33_ASAP7_75t_R n_9066 (.A1(n_8880_o_0),
    .A2(n_9062_o_0),
    .A3(n_9065_o_0),
    .B(n_8992_o_0),
    .Y(n_9066_o_0));
 OAI21xp33_ASAP7_75t_R n_9067 (.A1(n_9053_o_0),
    .A2(n_9059_o_0),
    .B(n_9066_o_0),
    .Y(n_9067_o_0));
 AOI21xp33_ASAP7_75t_R n_9068 (.A1(n_9048_o_0),
    .A2(n_9067_o_0),
    .B(n_8873_o_0),
    .Y(n_9068_o_0));
 AOI21xp33_ASAP7_75t_R n_9069 (.A1(n_8873_o_0),
    .A2(n_9025_o_0),
    .B(n_9068_o_0),
    .Y(n_9069_o_0));
 NOR2xp33_ASAP7_75t_R n_907 (.A(n_847_o_0),
    .B(n_836_o_0),
    .Y(n_907_o_0));
 NAND3xp33_ASAP7_75t_R n_9070 (.A(n_8945_o_0),
    .B(n_9018_o_0),
    .C(n_8942_o_0),
    .Y(n_9070_o_0));
 OAI31xp33_ASAP7_75t_R n_9071 (.A1(n_8939_o_0),
    .A2(n_9039_o_0),
    .A3(n_9041_o_0),
    .B(n_9070_o_0),
    .Y(n_9071_o_0));
 OAI21xp33_ASAP7_75t_R n_9072 (.A1(n_8943_o_0),
    .A2(n_8944_o_0),
    .B(n_8947_o_0),
    .Y(n_9072_o_0));
 INVx1_ASAP7_75t_R n_9073 (.A(n_9072_o_0),
    .Y(n_9073_o_0));
 OAI21xp33_ASAP7_75t_R n_9074 (.A1(n_8998_o_0),
    .A2(n_9073_o_0),
    .B(net64),
    .Y(n_9074_o_0));
 NOR2xp33_ASAP7_75t_R n_9075 (.A(n_8944_o_0),
    .B(n_9063_o_0),
    .Y(n_9075_o_0));
 OAI22xp33_ASAP7_75t_R n_9076 (.A1(n_9071_o_0),
    .A2(n_8889_o_0),
    .B1(n_9074_o_0),
    .B2(n_9075_o_0),
    .Y(n_9076_o_0));
 NAND2xp33_ASAP7_75t_R n_9077 (.A(n_8915_o_0),
    .B(n_8974_o_0),
    .Y(n_9077_o_0));
 INVx1_ASAP7_75t_R n_9078 (.A(n_9077_o_0),
    .Y(n_9078_o_0));
 OAI21xp33_ASAP7_75t_R n_9079 (.A1(n_8947_o_0),
    .A2(n_9078_o_0),
    .B(n_8964_o_0),
    .Y(n_9079_o_0));
 NOR2xp33_ASAP7_75t_R n_908 (.A(n_878_o_0),
    .B(n_907_o_0),
    .Y(n_908_o_0));
 AOI31xp33_ASAP7_75t_R n_9080 (.A1(n_8947_o_0),
    .A2(n_9012_o_0),
    .A3(n_8963_o_0),
    .B(n_8889_o_0),
    .Y(n_9080_o_0));
 OAI21xp33_ASAP7_75t_R n_9081 (.A1(n_8947_o_0),
    .A2(n_8974_o_0),
    .B(n_8968_o_0),
    .Y(n_9081_o_0));
 NOR2xp33_ASAP7_75t_R n_9082 (.A(net19),
    .B(n_8926_o_0),
    .Y(n_9082_o_0));
 AOI21xp33_ASAP7_75t_R n_9083 (.A1(n_8939_o_0),
    .A2(n_9082_o_0),
    .B(net64),
    .Y(n_9083_o_0));
 AOI21xp33_ASAP7_75t_R n_9084 (.A1(n_9081_o_0),
    .A2(n_9083_o_0),
    .B(n_8984_o_0),
    .Y(n_9084_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9085 (.A1(n_9044_o_0),
    .A2(n_9079_o_0),
    .B(n_9080_o_0),
    .C(n_9084_o_0),
    .D(n_9046_o_0),
    .Y(n_9085_o_0));
 OAI211xp5_ASAP7_75t_R n_9086 (.A1(n_8960_o_0),
    .A2(n_8947_o_0),
    .B(n_9004_o_0),
    .C(n_8942_o_0),
    .Y(n_9086_o_0));
 OAI31xp33_ASAP7_75t_R n_9087 (.A1(n_8939_o_0),
    .A2(n_8947_o_0),
    .A3(n_9029_o_0),
    .B(n_9086_o_0),
    .Y(n_9087_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9088 (.A1(n_8974_o_0),
    .A2(n_8915_o_0),
    .B(n_8926_o_0),
    .C(n_8939_o_0),
    .Y(n_9088_o_0));
 AOI21xp33_ASAP7_75t_R n_9089 (.A1(n_8915_o_0),
    .A2(n_8974_o_0),
    .B(n_8939_o_0),
    .Y(n_9089_o_0));
 HAxp5_ASAP7_75t_R n_909 (.A(n_859_o_0),
    .B(n_847_o_0),
    .CON(n_909_o_0),
    .SN(n_909_o_1));
 AOI21xp33_ASAP7_75t_R n_9090 (.A1(n_8926_o_0),
    .A2(n_9089_o_0),
    .B(n_8889_o_0),
    .Y(n_9090_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9091 (.A1(n_9088_o_0),
    .A2(n_8978_o_0),
    .B(n_9090_o_0),
    .C(n_8983_o_0),
    .Y(n_9091_o_0));
 OAI21xp33_ASAP7_75t_R n_9092 (.A1(n_9010_o_0),
    .A2(n_9087_o_0),
    .B(n_9091_o_0),
    .Y(n_9092_o_0));
 NOR2xp33_ASAP7_75t_R n_9093 (.A(n_8926_o_0),
    .B(n_8968_o_0),
    .Y(n_9093_o_0));
 INVx1_ASAP7_75t_R n_9094 (.A(n_9093_o_0),
    .Y(n_9094_o_0));
 OAI211xp5_ASAP7_75t_R n_9095 (.A1(net19),
    .A2(n_8947_o_0),
    .B(n_8995_o_0),
    .C(n_8963_o_0),
    .Y(n_9095_o_0));
 OAI21xp33_ASAP7_75t_R n_9096 (.A1(n_9012_o_0),
    .A2(n_9094_o_0),
    .B(n_9095_o_0),
    .Y(n_9096_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9097 (.A1(n_8915_o_0),
    .A2(net48),
    .B(n_8926_o_0),
    .C(n_8939_o_0),
    .Y(n_9097_o_0));
 AOI21xp33_ASAP7_75t_R n_9098 (.A1(n_9040_o_0),
    .A2(n_9097_o_0),
    .B(n_8889_o_0),
    .Y(n_9098_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9099 (.A1(n_9015_o_0),
    .A2(n_8970_o_0),
    .B(n_9098_o_0),
    .C(n_8880_o_0),
    .Y(n_9099_o_0));
 INVx1_ASAP7_75t_R n_910 (.A(n_907_o_0),
    .Y(n_910_o_0));
 OAI21xp33_ASAP7_75t_R n_9100 (.A1(n_9010_o_0),
    .A2(n_9096_o_0),
    .B(n_9099_o_0),
    .Y(n_9100_o_0));
 AOI21xp33_ASAP7_75t_R n_9101 (.A1(n_9092_o_0),
    .A2(n_9100_o_0),
    .B(n_8992_o_0),
    .Y(n_9101_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9102 (.A1(n_9008_o_0),
    .A2(n_9076_o_0),
    .B(n_9085_o_0),
    .C(n_9101_o_0),
    .Y(n_9102_o_0));
 NAND2xp33_ASAP7_75t_R n_9103 (.A(_00939_),
    .B(n_8871_o_0),
    .Y(n_9103_o_0));
 OAI21xp33_ASAP7_75t_R n_9104 (.A1(_00939_),
    .A2(n_8871_o_0),
    .B(n_9103_o_0),
    .Y(n_9104_o_0));
 INVx1_ASAP7_75t_R n_9105 (.A(n_9104_o_0),
    .Y(n_9105_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9106 (.A1(n_8974_o_0),
    .A2(n_8915_o_0),
    .B(n_8947_o_0),
    .C(n_8963_o_0),
    .Y(n_9106_o_0));
 AND3x1_ASAP7_75t_R n_9107 (.A(n_9086_o_0),
    .B(n_9037_o_0),
    .C(n_8992_o_0),
    .Y(n_9107_o_0));
 OAI31xp33_ASAP7_75t_R n_9108 (.A1(n_8939_o_0),
    .A2(n_8969_o_0),
    .A3(n_8970_o_0),
    .B(n_9015_o_0),
    .Y(n_9108_o_0));
 NOR3xp33_ASAP7_75t_R n_9109 (.A(n_9108_o_0),
    .B(n_9010_o_0),
    .C(n_8993_o_0),
    .Y(n_9109_o_0));
 AOI21xp33_ASAP7_75t_R n_911 (.A1(n_909_o_0),
    .A2(n_910_o_0),
    .B(n_877_o_0),
    .Y(n_911_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9110 (.A1(n_9060_o_0),
    .A2(n_9106_o_0),
    .B(n_9107_o_0),
    .C(n_9109_o_0),
    .Y(n_9110_o_0));
 AOI21xp33_ASAP7_75t_R n_9111 (.A1(n_8947_o_0),
    .A2(net19),
    .B(n_9013_o_0),
    .Y(n_9111_o_0));
 NOR2xp33_ASAP7_75t_R n_9112 (.A(n_8998_o_0),
    .B(n_9002_o_0),
    .Y(n_9112_o_0));
 AOI31xp33_ASAP7_75t_R n_9113 (.A1(n_8954_o_0),
    .A2(n_8958_o_0),
    .A3(n_8947_o_0),
    .B(n_8968_o_0),
    .Y(n_9113_o_0));
 AOI221xp5_ASAP7_75t_R n_9114 (.A1(n_8939_o_0),
    .A2(n_9039_o_0),
    .B1(n_9055_o_0),
    .B2(n_9054_o_0),
    .C(n_8972_o_0),
    .Y(n_9114_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9115 (.A1(n_8963_o_0),
    .A2(n_9040_o_0),
    .B(n_9113_o_0),
    .C(n_9114_o_0),
    .Y(n_9115_o_0));
 OAI31xp33_ASAP7_75t_R n_9116 (.A1(n_9037_o_0),
    .A2(n_9111_o_0),
    .A3(n_9112_o_0),
    .B(n_9115_o_0),
    .Y(n_9116_o_0));
 NAND2xp33_ASAP7_75t_R n_9117 (.A(n_8993_o_0),
    .B(n_9116_o_0),
    .Y(n_9117_o_0));
 AOI31xp33_ASAP7_75t_R n_9118 (.A1(n_8984_o_0),
    .A2(n_9110_o_0),
    .A3(n_9117_o_0),
    .B(n_8872_o_0),
    .Y(n_9118_o_0));
 NOR2xp33_ASAP7_75t_R n_9119 (.A(n_8952_o_0),
    .B(n_8998_o_0),
    .Y(n_9119_o_0));
 AOI211xp5_ASAP7_75t_R n_912 (.A1(n_908_o_0),
    .A2(n_909_o_0),
    .B(n_911_o_0),
    .C(net15),
    .Y(n_912_o_0));
 OAI31xp33_ASAP7_75t_R n_9120 (.A1(n_8926_o_0),
    .A2(n_8915_o_0),
    .A3(n_8904_o_0),
    .B(n_8942_o_0),
    .Y(n_9120_o_0));
 AOI21xp33_ASAP7_75t_R n_9121 (.A1(n_8948_o_0),
    .A2(n_9017_o_0),
    .B(n_9024_o_0),
    .Y(n_9121_o_0));
 OAI21xp33_ASAP7_75t_R n_9122 (.A1(n_8969_o_0),
    .A2(n_9120_o_0),
    .B(n_9121_o_0),
    .Y(n_9122_o_0));
 OAI31xp33_ASAP7_75t_R n_9123 (.A1(n_9046_o_0),
    .A2(n_9111_o_0),
    .A3(n_9119_o_0),
    .B(n_9122_o_0),
    .Y(n_9123_o_0));
 NAND2xp33_ASAP7_75t_R n_9124 (.A(net48),
    .B(n_8947_o_0),
    .Y(n_9124_o_0));
 OAI31xp33_ASAP7_75t_R n_9125 (.A1(n_8947_o_0),
    .A2(n_8946_o_0),
    .A3(n_8904_o_0),
    .B(n_8963_o_0),
    .Y(n_9125_o_0));
 OAI21xp33_ASAP7_75t_R n_9126 (.A1(n_9125_o_0),
    .A2(n_9049_o_0),
    .B(net64),
    .Y(n_9126_o_0));
 AOI31xp33_ASAP7_75t_R n_9127 (.A1(n_8942_o_0),
    .A2(n_9024_o_0),
    .A3(n_9124_o_0),
    .B(n_9126_o_0),
    .Y(n_9127_o_0));
 AOI211xp5_ASAP7_75t_R n_9128 (.A1(n_9123_o_0),
    .A2(n_9037_o_0),
    .B(n_8880_o_0),
    .C(n_9127_o_0),
    .Y(n_9128_o_0));
 INVx1_ASAP7_75t_R n_9129 (.A(n_9128_o_0),
    .Y(n_9129_o_0));
 NOR2xp67_ASAP7_75t_R n_913 (.A(n_847_o_0),
    .B(n_859_o_0),
    .Y(n_913_o_0));
 AOI22xp33_ASAP7_75t_R n_9130 (.A1(n_9102_o_0),
    .A2(n_9105_o_0),
    .B1(n_9118_o_0),
    .B2(n_9129_o_0),
    .Y(n_9130_o_0));
 NOR2xp33_ASAP7_75t_R n_9131 (.A(n_8904_o_0),
    .B(n_8947_o_0),
    .Y(n_9131_o_0));
 NAND2xp33_ASAP7_75t_R n_9132 (.A(net48),
    .B(n_8915_o_0),
    .Y(n_9132_o_0));
 INVx1_ASAP7_75t_R n_9133 (.A(n_9132_o_0),
    .Y(n_9133_o_0));
 OAI21xp33_ASAP7_75t_R n_9134 (.A1(n_9133_o_0),
    .A2(n_8947_o_0),
    .B(n_9113_o_0),
    .Y(n_9134_o_0));
 OAI31xp33_ASAP7_75t_R n_9135 (.A1(n_8939_o_0),
    .A2(n_9131_o_0),
    .A3(n_9060_o_0),
    .B(n_9134_o_0),
    .Y(n_9135_o_0));
 INVx1_ASAP7_75t_R n_9136 (.A(n_9064_o_0),
    .Y(n_9136_o_0));
 AOI21xp33_ASAP7_75t_R n_9137 (.A1(n_8947_o_0),
    .A2(net19),
    .B(n_9063_o_0),
    .Y(n_9137_o_0));
 OAI31xp33_ASAP7_75t_R n_9138 (.A1(n_8992_o_0),
    .A2(n_9136_o_0),
    .A3(n_9137_o_0),
    .B(n_9037_o_0),
    .Y(n_9138_o_0));
 AOI21xp33_ASAP7_75t_R n_9139 (.A1(n_9024_o_0),
    .A2(n_9135_o_0),
    .B(n_9138_o_0),
    .Y(n_9139_o_0));
 NAND2xp33_ASAP7_75t_R n_914 (.A(net32),
    .B(n_913_o_0),
    .Y(n_914_o_0));
 NOR2xp33_ASAP7_75t_R n_9140 (.A(n_8915_o_0),
    .B(n_8974_o_0),
    .Y(n_9140_o_0));
 NOR3xp33_ASAP7_75t_R n_9141 (.A(n_9140_o_0),
    .B(n_9131_o_0),
    .C(n_8968_o_0),
    .Y(n_9141_o_0));
 AOI211xp5_ASAP7_75t_R n_9142 (.A1(n_9124_o_0),
    .A2(n_8968_o_0),
    .B(n_9141_o_0),
    .C(n_9046_o_0),
    .Y(n_9142_o_0));
 OAI31xp33_ASAP7_75t_R n_9143 (.A1(net19),
    .A2(n_8947_o_0),
    .A3(n_8942_o_0),
    .B(n_8993_o_0),
    .Y(n_9143_o_0));
 AOI21xp33_ASAP7_75t_R n_9144 (.A1(n_9043_o_0),
    .A2(n_8964_o_0),
    .B(n_9143_o_0),
    .Y(n_9144_o_0));
 NOR3xp33_ASAP7_75t_R n_9145 (.A(n_9142_o_0),
    .B(n_9144_o_0),
    .C(n_9010_o_0),
    .Y(n_9145_o_0));
 NOR2xp33_ASAP7_75t_R n_9146 (.A(n_8926_o_0),
    .B(n_9012_o_0),
    .Y(n_9146_o_0));
 OAI21xp33_ASAP7_75t_R n_9147 (.A1(n_9146_o_0),
    .A2(n_9015_o_0),
    .B(n_9046_o_0),
    .Y(n_9147_o_0));
 NOR2xp33_ASAP7_75t_R n_9148 (.A(net19),
    .B(n_8947_o_0),
    .Y(n_9148_o_0));
 OAI22xp33_ASAP7_75t_R n_9149 (.A1(n_8976_o_0),
    .A2(n_8939_o_0),
    .B1(n_8968_o_0),
    .B2(n_9148_o_0),
    .Y(n_9149_o_0));
 NOR2xp33_ASAP7_75t_R n_915 (.A(n_881_o_0),
    .B(n_860_o_0),
    .Y(n_915_o_0));
 OAI22xp33_ASAP7_75t_R n_9150 (.A1(n_9147_o_0),
    .A2(n_8949_o_0),
    .B1(n_8993_o_0),
    .B2(n_9149_o_0),
    .Y(n_9150_o_0));
 OAI21xp33_ASAP7_75t_R n_9151 (.A1(n_9131_o_0),
    .A2(n_9120_o_0),
    .B(n_9024_o_0),
    .Y(n_9151_o_0));
 AO21x1_ASAP7_75t_R n_9152 (.A1(n_8968_o_0),
    .A2(n_9082_o_0),
    .B(n_9151_o_0),
    .Y(n_9152_o_0));
 AOI21xp33_ASAP7_75t_R n_9153 (.A1(n_8926_o_0),
    .A2(n_8915_o_0),
    .B(n_8968_o_0),
    .Y(n_9153_o_0));
 AOI21xp33_ASAP7_75t_R n_9154 (.A1(n_9153_o_0),
    .A2(n_9004_o_0),
    .B(n_9024_o_0),
    .Y(n_9154_o_0));
 OAI21xp33_ASAP7_75t_R n_9155 (.A1(n_9049_o_0),
    .A2(n_9125_o_0),
    .B(n_9154_o_0),
    .Y(n_9155_o_0));
 NAND3xp33_ASAP7_75t_R n_9156 (.A(n_9152_o_0),
    .B(n_9155_o_0),
    .C(n_9037_o_0),
    .Y(n_9156_o_0));
 OAI211xp5_ASAP7_75t_R n_9157 (.A1(n_9037_o_0),
    .A2(n_9150_o_0),
    .B(n_9156_o_0),
    .C(n_8983_o_0),
    .Y(n_9157_o_0));
 OAI31xp33_ASAP7_75t_R n_9158 (.A1(n_8983_o_0),
    .A2(n_9139_o_0),
    .A3(n_9145_o_0),
    .B(n_9157_o_0),
    .Y(n_9158_o_0));
 INVx1_ASAP7_75t_R n_9159 (.A(n_8994_o_0),
    .Y(n_9159_o_0));
 INVx1_ASAP7_75t_R n_916 (.A(n_915_o_0),
    .Y(n_916_o_0));
 OAI31xp33_ASAP7_75t_R n_9160 (.A1(n_8946_o_0),
    .A2(net19),
    .A3(n_8926_o_0),
    .B(n_8968_o_0),
    .Y(n_9160_o_0));
 NAND2xp33_ASAP7_75t_R n_9161 (.A(n_8904_o_0),
    .B(n_8947_o_0),
    .Y(n_9161_o_0));
 NAND3xp33_ASAP7_75t_R n_9162 (.A(n_9001_o_0),
    .B(n_9161_o_0),
    .C(n_8942_o_0),
    .Y(n_9162_o_0));
 OA211x2_ASAP7_75t_R n_9163 (.A1(n_9159_o_0),
    .A2(n_9160_o_0),
    .B(n_9162_o_0),
    .C(n_9037_o_0),
    .Y(n_9163_o_0));
 INVx1_ASAP7_75t_R n_9164 (.A(n_9113_o_0),
    .Y(n_9164_o_0));
 OAI21xp33_ASAP7_75t_R n_9165 (.A1(n_8946_o_0),
    .A2(n_8974_o_0),
    .B(n_8947_o_0),
    .Y(n_9165_o_0));
 NAND2xp33_ASAP7_75t_R n_9166 (.A(n_9165_o_0),
    .B(n_9017_o_0),
    .Y(n_9166_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9167 (.A1(n_9006_o_0),
    .A2(n_9164_o_0),
    .B(n_9166_o_0),
    .C(n_9010_o_0),
    .Y(n_9167_o_0));
 OR2x2_ASAP7_75t_R n_9168 (.A(n_8924_o_0),
    .B(n_8923_o_0),
    .Y(n_9168_o_0));
 AOI211xp5_ASAP7_75t_R n_9169 (.A1(n_8925_o_0),
    .A2(n_9168_o_0),
    .B(n_8974_o_0),
    .C(n_8946_o_0),
    .Y(n_9169_o_0));
 NOR2xp33_ASAP7_75t_R n_917 (.A(n_847_o_0),
    .B(n_864_o_0),
    .Y(n_917_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9170 (.A1(n_9160_o_0),
    .A2(n_9169_o_0),
    .B(n_9037_o_0),
    .C(n_9046_o_0),
    .Y(n_9170_o_0));
 NAND3xp33_ASAP7_75t_R n_9171 (.A(n_9018_o_0),
    .B(n_8994_o_0),
    .C(n_8942_o_0),
    .Y(n_9171_o_0));
 NOR4xp25_ASAP7_75t_R n_9172 (.A(n_9159_o_0),
    .B(n_9046_o_0),
    .C(n_8976_o_0),
    .D(n_8968_o_0),
    .Y(n_9172_o_0));
 AOI211xp5_ASAP7_75t_R n_9173 (.A1(n_8915_o_0),
    .A2(n_8947_o_0),
    .B(n_8963_o_0),
    .C(net19),
    .Y(n_9173_o_0));
 OAI21xp33_ASAP7_75t_R n_9174 (.A1(n_9173_o_0),
    .A2(n_9026_o_0),
    .B(n_8972_o_0),
    .Y(n_9174_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9175 (.A1(n_9170_o_0),
    .A2(n_9171_o_0),
    .B(n_9172_o_0),
    .C(n_9174_o_0),
    .Y(n_9175_o_0));
 OAI31xp33_ASAP7_75t_R n_9176 (.A1(n_8992_o_0),
    .A2(n_9163_o_0),
    .A3(n_9167_o_0),
    .B(n_9175_o_0),
    .Y(n_9176_o_0));
 OA21x2_ASAP7_75t_R n_9177 (.A1(n_9176_o_0),
    .A2(n_9008_o_0),
    .B(n_9104_o_0),
    .Y(n_9177_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9178 (.A1(n_8947_o_0),
    .A2(n_9012_o_0),
    .B(n_9013_o_0),
    .C(n_8889_o_0),
    .Y(n_9178_o_0));
 NOR2xp33_ASAP7_75t_R n_9179 (.A(n_9131_o_0),
    .B(n_9120_o_0),
    .Y(n_9179_o_0));
 INVx1_ASAP7_75t_R n_918 (.A(n_917_o_0),
    .Y(n_918_o_0));
 AOI211xp5_ASAP7_75t_R n_9180 (.A1(n_9029_o_0),
    .A2(n_8926_o_0),
    .B(n_8939_o_0),
    .C(n_9016_o_0),
    .Y(n_9180_o_0));
 OAI21xp33_ASAP7_75t_R n_9181 (.A1(n_9179_o_0),
    .A2(n_9180_o_0),
    .B(n_9037_o_0),
    .Y(n_9181_o_0));
 OAI21xp33_ASAP7_75t_R n_9182 (.A1(n_9136_o_0),
    .A2(n_9178_o_0),
    .B(n_9181_o_0),
    .Y(n_9182_o_0));
 NAND2xp33_ASAP7_75t_R n_9183 (.A(n_9161_o_0),
    .B(n_8959_o_0),
    .Y(n_9183_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9184 (.A1(n_8968_o_0),
    .A2(n_9159_o_0),
    .B(n_9183_o_0),
    .C(n_9002_o_0),
    .Y(n_9184_o_0));
 INVx1_ASAP7_75t_R n_9185 (.A(n_8979_o_0),
    .Y(n_9185_o_0));
 NOR3xp33_ASAP7_75t_R n_9186 (.A(n_9005_o_0),
    .B(n_9185_o_0),
    .C(n_8968_o_0),
    .Y(n_9186_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9187 (.A1(n_8963_o_0),
    .A2(n_9018_o_0),
    .B(n_9186_o_0),
    .C(n_8889_o_0),
    .Y(n_9187_o_0));
 OAI211xp5_ASAP7_75t_R n_9188 (.A1(n_8889_o_0),
    .A2(n_9184_o_0),
    .B(n_9187_o_0),
    .C(n_8993_o_0),
    .Y(n_9188_o_0));
 OAI211xp5_ASAP7_75t_R n_9189 (.A1(n_9182_o_0),
    .A2(n_9046_o_0),
    .B(n_9188_o_0),
    .C(n_8983_o_0),
    .Y(n_9189_o_0));
 NAND2xp33_ASAP7_75t_R n_919 (.A(n_881_o_0),
    .B(n_918_o_0),
    .Y(n_919_o_0));
 AOI22xp33_ASAP7_75t_R n_9190 (.A1(n_9158_o_0),
    .A2(n_8872_o_0),
    .B1(n_9177_o_0),
    .B2(n_9189_o_0),
    .Y(n_9190_o_0));
 OAI21xp33_ASAP7_75t_R n_9191 (.A1(n_8963_o_0),
    .A2(n_9001_o_0),
    .B(n_8993_o_0),
    .Y(n_9191_o_0));
 OAI21xp33_ASAP7_75t_R n_9192 (.A1(net48),
    .A2(n_8946_o_0),
    .B(n_8947_o_0),
    .Y(n_9192_o_0));
 AOI21xp33_ASAP7_75t_R n_9193 (.A1(n_9192_o_0),
    .A2(n_9153_o_0),
    .B(n_8993_o_0),
    .Y(n_9193_o_0));
 OAI31xp33_ASAP7_75t_R n_9194 (.A1(n_8939_o_0),
    .A2(n_9006_o_0),
    .A3(n_8970_o_0),
    .B(n_9193_o_0),
    .Y(n_9194_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9195 (.A1(n_9017_o_0),
    .A2(n_9165_o_0),
    .B(n_9191_o_0),
    .C(n_9194_o_0),
    .Y(n_9195_o_0));
 OAI21xp33_ASAP7_75t_R n_9196 (.A1(n_8942_o_0),
    .A2(n_8945_o_0),
    .B(n_8993_o_0),
    .Y(n_9196_o_0));
 NOR2xp33_ASAP7_75t_R n_9197 (.A(net19),
    .B(n_8947_o_0),
    .Y(n_9197_o_0));
 AOI31xp33_ASAP7_75t_R n_9198 (.A1(n_8939_o_0),
    .A2(n_8960_o_0),
    .A3(n_8947_o_0),
    .B(n_9046_o_0),
    .Y(n_9198_o_0));
 OAI31xp33_ASAP7_75t_R n_9199 (.A1(n_8939_o_0),
    .A2(n_9197_o_0),
    .A3(n_9049_o_0),
    .B(n_9198_o_0),
    .Y(n_9199_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_920 (.A1(n_916_o_0),
    .A2(n_919_o_0),
    .B(n_877_o_0),
    .C(n_891_o_0),
    .Y(n_920_o_0));
 AOI21xp33_ASAP7_75t_R n_9200 (.A1(n_9196_o_0),
    .A2(n_9199_o_0),
    .B(n_9052_o_0),
    .Y(n_9200_o_0));
 AOI21xp33_ASAP7_75t_R n_9201 (.A1(n_8889_o_0),
    .A2(n_9195_o_0),
    .B(n_9200_o_0),
    .Y(n_9201_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9202 (.A1(n_8926_o_0),
    .A2(n_8960_o_0),
    .B(n_8942_o_0),
    .C(n_9078_o_0),
    .Y(n_9202_o_0));
 OAI31xp33_ASAP7_75t_R n_9203 (.A1(n_8947_o_0),
    .A2(n_8960_o_0),
    .A3(n_8942_o_0),
    .B(n_9077_o_0),
    .Y(n_9203_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9204 (.A1(n_8926_o_0),
    .A2(n_8915_o_0),
    .B(n_9001_o_0),
    .C(n_8963_o_0),
    .Y(n_9204_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9205 (.A1(n_9202_o_0),
    .A2(n_9203_o_0),
    .B(n_9204_o_0),
    .C(n_9037_o_0),
    .Y(n_9205_o_0));
 AO21x1_ASAP7_75t_R n_9206 (.A1(n_9095_o_0),
    .A2(n_9042_o_0),
    .B(n_9037_o_0),
    .Y(n_9206_o_0));
 AOI21xp33_ASAP7_75t_R n_9207 (.A1(n_9165_o_0),
    .A2(n_9153_o_0),
    .B(n_9010_o_0),
    .Y(n_9207_o_0));
 OAI21xp33_ASAP7_75t_R n_9208 (.A1(n_9049_o_0),
    .A2(n_9125_o_0),
    .B(n_9207_o_0),
    .Y(n_9208_o_0));
 OAI31xp33_ASAP7_75t_R n_9209 (.A1(n_9160_o_0),
    .A2(n_9159_o_0),
    .A3(n_8972_o_0),
    .B(n_9208_o_0),
    .Y(n_9209_o_0));
 AOI31xp33_ASAP7_75t_R n_921 (.A1(n_877_o_0),
    .A2(n_914_o_0),
    .A3(n_882_o_0),
    .B(n_920_o_0),
    .Y(n_921_o_0));
 AOI321xp33_ASAP7_75t_R n_9210 (.A1(n_9205_o_0),
    .A2(n_9206_o_0),
    .A3(n_8993_o_0),
    .B1(n_9024_o_0),
    .B2(n_9209_o_0),
    .C(n_9008_o_0),
    .Y(n_9210_o_0));
 AOI21xp33_ASAP7_75t_R n_9211 (.A1(n_8983_o_0),
    .A2(n_9201_o_0),
    .B(n_9210_o_0),
    .Y(n_9211_o_0));
 AO21x1_ASAP7_75t_R n_9212 (.A1(n_8960_o_0),
    .A2(n_8947_o_0),
    .B(n_9125_o_0),
    .Y(n_9212_o_0));
 OAI31xp33_ASAP7_75t_R n_9213 (.A1(n_8968_o_0),
    .A2(n_8976_o_0),
    .A3(n_9169_o_0),
    .B(n_9212_o_0),
    .Y(n_9213_o_0));
 AOI21xp33_ASAP7_75t_R n_9214 (.A1(n_8926_o_0),
    .A2(n_8960_o_0),
    .B(n_8942_o_0),
    .Y(n_9214_o_0));
 AOI211xp5_ASAP7_75t_R n_9215 (.A1(n_9214_o_0),
    .A2(n_8928_o_0),
    .B(n_8972_o_0),
    .C(n_8996_o_0),
    .Y(n_9215_o_0));
 AOI21xp33_ASAP7_75t_R n_9216 (.A1(n_8889_o_0),
    .A2(n_9213_o_0),
    .B(n_9215_o_0),
    .Y(n_9216_o_0));
 AOI21xp33_ASAP7_75t_R n_9217 (.A1(n_9165_o_0),
    .A2(n_8959_o_0),
    .B(n_8889_o_0),
    .Y(n_9217_o_0));
 OAI21xp33_ASAP7_75t_R n_9218 (.A1(n_9088_o_0),
    .A2(n_8978_o_0),
    .B(n_9217_o_0),
    .Y(n_9218_o_0));
 OAI21xp33_ASAP7_75t_R n_9219 (.A1(n_9140_o_0),
    .A2(n_9041_o_0),
    .B(n_8968_o_0),
    .Y(n_9219_o_0));
 OAI21xp33_ASAP7_75t_R n_922 (.A1(n_912_o_0),
    .A2(n_921_o_0),
    .B(n_904_o_0),
    .Y(n_922_o_0));
 NAND3xp33_ASAP7_75t_R n_9220 (.A(n_9219_o_0),
    .B(n_9120_o_0),
    .C(net64),
    .Y(n_9220_o_0));
 AOI21xp33_ASAP7_75t_R n_9221 (.A1(n_9218_o_0),
    .A2(n_9220_o_0),
    .B(n_8993_o_0),
    .Y(n_9221_o_0));
 AOI211xp5_ASAP7_75t_R n_9222 (.A1(n_9046_o_0),
    .A2(n_9216_o_0),
    .B(n_9221_o_0),
    .C(n_8983_o_0),
    .Y(n_9222_o_0));
 OAI31xp33_ASAP7_75t_R n_9223 (.A1(n_8968_o_0),
    .A2(n_9185_o_0),
    .A3(n_9146_o_0),
    .B(n_9183_o_0),
    .Y(n_9223_o_0));
 NAND3xp33_ASAP7_75t_R n_9224 (.A(n_8945_o_0),
    .B(n_9161_o_0),
    .C(n_8942_o_0),
    .Y(n_9224_o_0));
 AOI21xp33_ASAP7_75t_R n_9225 (.A1(n_9219_o_0),
    .A2(n_9224_o_0),
    .B(n_8993_o_0),
    .Y(n_9225_o_0));
 AOI21xp33_ASAP7_75t_R n_9226 (.A1(n_8993_o_0),
    .A2(n_9223_o_0),
    .B(n_9225_o_0),
    .Y(n_9226_o_0));
 AOI31xp33_ASAP7_75t_R n_9227 (.A1(n_8939_o_0),
    .A2(n_8958_o_0),
    .A3(n_8954_o_0),
    .B(n_8926_o_0),
    .Y(n_9227_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9228 (.A1(n_8963_o_0),
    .A2(n_9051_o_0),
    .B(n_8926_o_0),
    .C(n_9227_o_0),
    .Y(n_9228_o_0));
 OAI21xp33_ASAP7_75t_R n_9229 (.A1(n_8946_o_0),
    .A2(n_8926_o_0),
    .B(n_8968_o_0),
    .Y(n_9229_o_0));
 INVx1_ASAP7_75t_R n_923 (.A(_00978_),
    .Y(n_923_o_0));
 AOI21xp33_ASAP7_75t_R n_9230 (.A1(n_9132_o_0),
    .A2(n_8926_o_0),
    .B(n_9229_o_0),
    .Y(n_9230_o_0));
 OAI221xp5_ASAP7_75t_R n_9231 (.A1(n_8952_o_0),
    .A2(n_8998_o_0),
    .B1(n_8963_o_0),
    .B2(n_9072_o_0),
    .C(n_9024_o_0),
    .Y(n_9231_o_0));
 OAI31xp33_ASAP7_75t_R n_9232 (.A1(n_8992_o_0),
    .A2(n_9228_o_0),
    .A3(n_9230_o_0),
    .B(n_9231_o_0),
    .Y(n_9232_o_0));
 OAI22xp33_ASAP7_75t_R n_9233 (.A1(n_9232_o_0),
    .A2(n_8889_o_0),
    .B1(n_8879_o_0),
    .B2(n_8878_o_0),
    .Y(n_9233_o_0));
 AOI21xp33_ASAP7_75t_R n_9234 (.A1(net64),
    .A2(n_9226_o_0),
    .B(n_9233_o_0),
    .Y(n_9234_o_0));
 OAI21xp33_ASAP7_75t_R n_9235 (.A1(n_9222_o_0),
    .A2(n_9234_o_0),
    .B(n_8872_o_0),
    .Y(n_9235_o_0));
 OAI21xp33_ASAP7_75t_R n_9236 (.A1(n_9105_o_0),
    .A2(n_9211_o_0),
    .B(n_9235_o_0),
    .Y(n_9236_o_0));
 AO21x1_ASAP7_75t_R n_9237 (.A1(net19),
    .A2(n_8926_o_0),
    .B(n_9057_o_0),
    .Y(n_9237_o_0));
 AOI21xp33_ASAP7_75t_R n_9238 (.A1(n_9055_o_0),
    .A2(n_9029_o_0),
    .B(net64),
    .Y(n_9238_o_0));
 NOR3xp33_ASAP7_75t_R n_9239 (.A(n_9113_o_0),
    .B(n_9010_o_0),
    .C(n_9089_o_0),
    .Y(n_9239_o_0));
 XNOR2xp5_ASAP7_75t_R n_924 (.A(_00444_),
    .B(_00882_),
    .Y(n_924_o_0));
 AOI21xp33_ASAP7_75t_R n_9240 (.A1(n_9237_o_0),
    .A2(n_9238_o_0),
    .B(n_9239_o_0),
    .Y(n_9240_o_0));
 INVx1_ASAP7_75t_R n_9241 (.A(n_9061_o_0),
    .Y(n_9241_o_0));
 AOI21xp33_ASAP7_75t_R n_9242 (.A1(n_8958_o_0),
    .A2(n_9033_o_0),
    .B(n_8939_o_0),
    .Y(n_9242_o_0));
 NOR2xp33_ASAP7_75t_R n_9243 (.A(n_8972_o_0),
    .B(n_9242_o_0),
    .Y(n_9243_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9244 (.A1(n_8915_o_0),
    .A2(n_8926_o_0),
    .B(n_9057_o_0),
    .C(n_9243_o_0),
    .Y(n_9244_o_0));
 OAI31xp33_ASAP7_75t_R n_9245 (.A1(n_9037_o_0),
    .A2(n_9241_o_0),
    .A3(n_8996_o_0),
    .B(n_9244_o_0),
    .Y(n_9245_o_0));
 OAI21xp33_ASAP7_75t_R n_9246 (.A1(n_8993_o_0),
    .A2(n_9245_o_0),
    .B(n_9008_o_0),
    .Y(n_9246_o_0));
 AOI21xp33_ASAP7_75t_R n_9247 (.A1(n_9046_o_0),
    .A2(n_9240_o_0),
    .B(n_9246_o_0),
    .Y(n_9247_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9248 (.A1(n_8947_o_0),
    .A2(n_9054_o_0),
    .B(n_9161_o_0),
    .C(n_8942_o_0),
    .Y(n_9248_o_0));
 OAI21xp33_ASAP7_75t_R n_9249 (.A1(n_9248_o_0),
    .A2(n_9111_o_0),
    .B(n_9037_o_0),
    .Y(n_9249_o_0));
 XNOR2xp5_ASAP7_75t_R n_925 (.A(_00914_),
    .B(n_924_o_0),
    .Y(n_925_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9250 (.A1(n_8999_o_0),
    .A2(n_9192_o_0),
    .B(n_9093_o_0),
    .C(n_8889_o_0),
    .Y(n_9250_o_0));
 OAI21xp33_ASAP7_75t_R n_9251 (.A1(n_8926_o_0),
    .A2(n_8960_o_0),
    .B(n_9097_o_0),
    .Y(n_9251_o_0));
 OAI31xp33_ASAP7_75t_R n_9252 (.A1(n_8968_o_0),
    .A2(n_8969_o_0),
    .A3(n_8970_o_0),
    .B(n_9251_o_0),
    .Y(n_9252_o_0));
 OAI21xp33_ASAP7_75t_R n_9253 (.A1(n_8926_o_0),
    .A2(n_9077_o_0),
    .B(n_8942_o_0),
    .Y(n_9253_o_0));
 OAI21xp33_ASAP7_75t_R n_9254 (.A1(n_8926_o_0),
    .A2(n_9054_o_0),
    .B(n_8968_o_0),
    .Y(n_9254_o_0));
 AOI21xp33_ASAP7_75t_R n_9255 (.A1(n_9253_o_0),
    .A2(n_9254_o_0),
    .B(n_8889_o_0),
    .Y(n_9255_o_0));
 AOI211xp5_ASAP7_75t_R n_9256 (.A1(n_8889_o_0),
    .A2(n_9252_o_0),
    .B(n_9255_o_0),
    .C(n_9024_o_0),
    .Y(n_9256_o_0));
 AOI31xp33_ASAP7_75t_R n_9257 (.A1(n_9024_o_0),
    .A2(n_9249_o_0),
    .A3(n_9250_o_0),
    .B(n_9256_o_0),
    .Y(n_9257_o_0));
 OAI21xp33_ASAP7_75t_R n_9258 (.A1(n_8983_o_0),
    .A2(n_9257_o_0),
    .B(n_8873_o_0),
    .Y(n_9258_o_0));
 AOI211xp5_ASAP7_75t_R n_9259 (.A1(n_8947_o_0),
    .A2(net19),
    .B(n_9056_o_0),
    .C(n_8963_o_0),
    .Y(n_9259_o_0));
 INVx1_ASAP7_75t_R n_926 (.A(n_925_o_0),
    .Y(n_926_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9260 (.A1(n_8952_o_0),
    .A2(n_9039_o_0),
    .B(n_8939_o_0),
    .C(n_9037_o_0),
    .Y(n_9260_o_0));
 NAND2xp33_ASAP7_75t_R n_9261 (.A(n_9260_o_0),
    .B(n_9044_o_0),
    .Y(n_9261_o_0));
 OAI31xp33_ASAP7_75t_R n_9262 (.A1(net64),
    .A2(n_9180_o_0),
    .A3(n_9259_o_0),
    .B(n_9261_o_0),
    .Y(n_9262_o_0));
 NOR2xp33_ASAP7_75t_R n_9263 (.A(n_9106_o_0),
    .B(n_9073_o_0),
    .Y(n_9263_o_0));
 NOR3xp33_ASAP7_75t_R n_9264 (.A(n_9132_o_0),
    .B(n_8947_o_0),
    .C(n_8972_o_0),
    .Y(n_9264_o_0));
 AOI211xp5_ASAP7_75t_R n_9265 (.A1(_00935_),
    .A2(n_8935_o_0),
    .B(n_8926_o_0),
    .C(n_8938_o_0),
    .Y(n_9265_o_0));
 AOI311xp33_ASAP7_75t_R n_9266 (.A1(n_8958_o_0),
    .A2(n_8954_o_0),
    .A3(n_9265_o_0),
    .B(n_8972_o_0),
    .C(n_9169_o_0),
    .Y(n_9266_o_0));
 OAI211xp5_ASAP7_75t_R n_9267 (.A1(n_9169_o_0),
    .A2(n_8976_o_0),
    .B(n_8968_o_0),
    .C(n_9046_o_0),
    .Y(n_9267_o_0));
 AOI31xp33_ASAP7_75t_R n_9268 (.A1(n_8958_o_0),
    .A2(n_9265_o_0),
    .A3(n_8954_o_0),
    .B(n_8972_o_0),
    .Y(n_9268_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9269 (.A1(n_8963_o_0),
    .A2(n_9001_o_0),
    .B(n_9268_o_0),
    .C(n_9046_o_0),
    .Y(n_9269_o_0));
 XNOR2xp5_ASAP7_75t_R n_927 (.A(_00946_),
    .B(n_926_o_0),
    .Y(n_927_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9270 (.A1(n_9264_o_0),
    .A2(n_8963_o_0),
    .B(n_9266_o_0),
    .C(n_9267_o_0),
    .D(n_9269_o_0),
    .Y(n_9270_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9271 (.A1(n_9058_o_0),
    .A2(n_9263_o_0),
    .B(n_9270_o_0),
    .C(n_8880_o_0),
    .Y(n_9271_o_0));
 OAI21xp33_ASAP7_75t_R n_9272 (.A1(n_8993_o_0),
    .A2(n_9262_o_0),
    .B(n_9271_o_0),
    .Y(n_9272_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9273 (.A1(n_8974_o_0),
    .A2(n_8947_o_0),
    .B(n_9063_o_0),
    .C(n_9121_o_0),
    .Y(n_9273_o_0));
 OAI31xp33_ASAP7_75t_R n_9274 (.A1(n_9046_o_0),
    .A2(n_9119_o_0),
    .A3(n_9141_o_0),
    .B(n_9273_o_0),
    .Y(n_9274_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9275 (.A1(n_8947_o_0),
    .A2(n_9051_o_0),
    .B(n_9057_o_0),
    .C(n_9024_o_0),
    .Y(n_9275_o_0));
 NOR2xp33_ASAP7_75t_R n_9276 (.A(n_9131_o_0),
    .B(n_9060_o_0),
    .Y(n_9276_o_0));
 AOI211xp5_ASAP7_75t_R n_9277 (.A1(n_9276_o_0),
    .A2(n_8939_o_0),
    .B(n_9046_o_0),
    .C(n_9242_o_0),
    .Y(n_9277_o_0));
 OAI21xp33_ASAP7_75t_R n_9278 (.A1(n_9275_o_0),
    .A2(n_9277_o_0),
    .B(n_9010_o_0),
    .Y(n_9278_o_0));
 OAI211xp5_ASAP7_75t_R n_9279 (.A1(n_9010_o_0),
    .A2(n_9274_o_0),
    .B(n_9278_o_0),
    .C(n_8984_o_0),
    .Y(n_9279_o_0));
 NOR2xp33_ASAP7_75t_R n_928 (.A(n_923_o_0),
    .B(n_927_o_0),
    .Y(n_928_o_0));
 NAND3xp33_ASAP7_75t_R n_9280 (.A(n_9272_o_0),
    .B(n_9279_o_0),
    .C(n_9105_o_0),
    .Y(n_9280_o_0));
 OAI21xp33_ASAP7_75t_R n_9281 (.A1(n_9247_o_0),
    .A2(n_9258_o_0),
    .B(n_9280_o_0),
    .Y(n_9281_o_0));
 AOI21xp33_ASAP7_75t_R n_9282 (.A1(n_8926_o_0),
    .A2(n_9077_o_0),
    .B(n_8963_o_0),
    .Y(n_9282_o_0));
 OAI21xp33_ASAP7_75t_R n_9283 (.A1(n_8944_o_0),
    .A2(n_9011_o_0),
    .B(n_9010_o_0),
    .Y(n_9283_o_0));
 AOI21xp33_ASAP7_75t_R n_9284 (.A1(n_8928_o_0),
    .A2(n_9282_o_0),
    .B(n_9283_o_0),
    .Y(n_9284_o_0));
 AOI211xp5_ASAP7_75t_R n_9285 (.A1(net19),
    .A2(n_8939_o_0),
    .B(n_9242_o_0),
    .C(n_9037_o_0),
    .Y(n_9285_o_0));
 OR3x1_ASAP7_75t_R n_9286 (.A(n_9284_o_0),
    .B(n_9285_o_0),
    .C(n_9024_o_0),
    .Y(n_9286_o_0));
 OAI32xp33_ASAP7_75t_R n_9287 (.A1(n_8963_o_0),
    .A2(n_8926_o_0),
    .A3(n_8960_o_0),
    .B1(n_9254_o_0),
    .B2(n_9197_o_0),
    .Y(n_9287_o_0));
 OAI21xp33_ASAP7_75t_R n_9288 (.A1(n_9060_o_0),
    .A2(n_9015_o_0),
    .B(n_9160_o_0),
    .Y(n_9288_o_0));
 OAI21xp33_ASAP7_75t_R n_9289 (.A1(n_9010_o_0),
    .A2(n_9288_o_0),
    .B(n_9024_o_0),
    .Y(n_9289_o_0));
 AOI211xp5_ASAP7_75t_R n_929 (.A1(n_923_o_0),
    .A2(n_927_o_0),
    .B(n_928_o_0),
    .C(ld),
    .Y(n_929_o_0));
 AO21x1_ASAP7_75t_R n_9290 (.A1(n_9037_o_0),
    .A2(n_9287_o_0),
    .B(n_9289_o_0),
    .Y(n_9290_o_0));
 OAI21xp33_ASAP7_75t_R n_9291 (.A1(n_9204_o_0),
    .A2(n_9214_o_0),
    .B(net64),
    .Y(n_9291_o_0));
 AO21x1_ASAP7_75t_R n_9292 (.A1(n_9029_o_0),
    .A2(n_8947_o_0),
    .B(n_9097_o_0),
    .Y(n_9292_o_0));
 AOI21xp33_ASAP7_75t_R n_9293 (.A1(n_9010_o_0),
    .A2(n_9292_o_0),
    .B(n_8993_o_0),
    .Y(n_9293_o_0));
 AOI211xp5_ASAP7_75t_R n_9294 (.A1(n_8947_o_0),
    .A2(net19),
    .B(n_8963_o_0),
    .C(n_8915_o_0),
    .Y(n_9294_o_0));
 NOR3xp33_ASAP7_75t_R n_9295 (.A(n_9056_o_0),
    .B(n_8942_o_0),
    .C(n_8927_o_0),
    .Y(n_9295_o_0));
 NOR2xp33_ASAP7_75t_R n_9296 (.A(n_9010_o_0),
    .B(n_8975_o_0),
    .Y(n_9296_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9297 (.A1(n_8926_o_0),
    .A2(n_9029_o_0),
    .B(n_9088_o_0),
    .C(n_9296_o_0),
    .Y(n_9297_o_0));
 OAI31xp33_ASAP7_75t_R n_9298 (.A1(net64),
    .A2(n_9294_o_0),
    .A3(n_9295_o_0),
    .B(n_9297_o_0),
    .Y(n_9298_o_0));
 AOI221xp5_ASAP7_75t_R n_9299 (.A1(n_9291_o_0),
    .A2(n_9293_o_0),
    .B1(n_8993_o_0),
    .B2(n_9298_o_0),
    .C(n_8983_o_0),
    .Y(n_9299_o_0));
 AOI21xp33_ASAP7_75t_R n_930 (.A1(key[22]),
    .A2(ld),
    .B(n_929_o_0),
    .Y(n_930_o_0));
 AOI31xp33_ASAP7_75t_R n_9300 (.A1(n_9008_o_0),
    .A2(n_9286_o_0),
    .A3(n_9290_o_0),
    .B(n_9299_o_0),
    .Y(n_9300_o_0));
 INVx1_ASAP7_75t_R n_9301 (.A(n_9125_o_0),
    .Y(n_9301_o_0));
 AOI21xp33_ASAP7_75t_R n_9302 (.A1(n_9018_o_0),
    .A2(n_9301_o_0),
    .B(n_9153_o_0),
    .Y(n_9302_o_0));
 AOI22xp33_ASAP7_75t_R n_9303 (.A1(n_9302_o_0),
    .A2(net64),
    .B1(n_9088_o_0),
    .B2(n_9080_o_0),
    .Y(n_9303_o_0));
 AOI21xp33_ASAP7_75t_R n_9304 (.A1(n_9132_o_0),
    .A2(n_8942_o_0),
    .B(n_9301_o_0),
    .Y(n_9304_o_0));
 OAI311xp33_ASAP7_75t_R n_9305 (.A1(n_8943_o_0),
    .A2(n_8944_o_0),
    .A3(n_8947_o_0),
    .B1(n_9192_o_0),
    .C1(n_8963_o_0),
    .Y(n_9305_o_0));
 OAI31xp33_ASAP7_75t_R n_9306 (.A1(n_8968_o_0),
    .A2(n_9006_o_0),
    .A3(n_9049_o_0),
    .B(n_9305_o_0),
    .Y(n_9306_o_0));
 AOI21xp33_ASAP7_75t_R n_9307 (.A1(n_9010_o_0),
    .A2(n_9306_o_0),
    .B(n_8993_o_0),
    .Y(n_9307_o_0));
 OAI21xp33_ASAP7_75t_R n_9308 (.A1(n_9037_o_0),
    .A2(n_9304_o_0),
    .B(n_9307_o_0),
    .Y(n_9308_o_0));
 OAI21xp33_ASAP7_75t_R n_9309 (.A1(n_9303_o_0),
    .A2(n_9024_o_0),
    .B(n_9308_o_0),
    .Y(n_9309_o_0));
 INVx1_ASAP7_75t_R n_931 (.A(n_930_o_0),
    .Y(n_931_o_0));
 AOI21xp33_ASAP7_75t_R n_9310 (.A1(n_8926_o_0),
    .A2(n_8960_o_0),
    .B(n_9120_o_0),
    .Y(n_9310_o_0));
 AOI31xp33_ASAP7_75t_R n_9311 (.A1(n_8963_o_0),
    .A2(n_8977_o_0),
    .A3(n_9165_o_0),
    .B(n_9310_o_0),
    .Y(n_9311_o_0));
 OAI21xp33_ASAP7_75t_R n_9312 (.A1(n_8998_o_0),
    .A2(n_9140_o_0),
    .B(n_8972_o_0),
    .Y(n_9312_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9313 (.A1(n_8942_o_0),
    .A2(n_8915_o_0),
    .B(n_9312_o_0),
    .C(n_8993_o_0),
    .Y(n_9313_o_0));
 AOI21xp33_ASAP7_75t_R n_9314 (.A1(n_9037_o_0),
    .A2(n_9311_o_0),
    .B(n_9313_o_0),
    .Y(n_9314_o_0));
 INVx1_ASAP7_75t_R n_9315 (.A(n_9017_o_0),
    .Y(n_9315_o_0));
 OAI21xp33_ASAP7_75t_R n_9316 (.A1(n_9125_o_0),
    .A2(n_9016_o_0),
    .B(n_9037_o_0),
    .Y(n_9316_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9317 (.A1(n_9132_o_0),
    .A2(n_9093_o_0),
    .B(n_9316_o_0),
    .C(n_9024_o_0),
    .Y(n_9317_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9318 (.A1(n_9315_o_0),
    .A2(n_9146_o_0),
    .B(n_9030_o_0),
    .C(n_9317_o_0),
    .Y(n_9318_o_0));
 OAI31xp33_ASAP7_75t_R n_9319 (.A1(n_9008_o_0),
    .A2(n_9314_o_0),
    .A3(n_9318_o_0),
    .B(n_9104_o_0),
    .Y(n_9319_o_0));
 AOI21xp33_ASAP7_75t_R n_932 (.A1(n_906_o_0),
    .A2(n_922_o_0),
    .B(n_931_o_0),
    .Y(n_932_o_0));
 AO21x1_ASAP7_75t_R n_9320 (.A1(n_9309_o_0),
    .A2(n_8983_o_0),
    .B(n_9319_o_0),
    .Y(n_9320_o_0));
 OAI21xp33_ASAP7_75t_R n_9321 (.A1(n_8873_o_0),
    .A2(n_9300_o_0),
    .B(n_9320_o_0),
    .Y(n_9321_o_0));
 OAI21xp33_ASAP7_75t_R n_9322 (.A1(n_8939_o_0),
    .A2(n_9049_o_0),
    .B(n_9237_o_0),
    .Y(n_9322_o_0));
 AOI21xp33_ASAP7_75t_R n_9323 (.A1(n_9010_o_0),
    .A2(n_9322_o_0),
    .B(n_8993_o_0),
    .Y(n_9323_o_0));
 AOI21xp33_ASAP7_75t_R n_9324 (.A1(net19),
    .A2(n_8926_o_0),
    .B(n_8939_o_0),
    .Y(n_9324_o_0));
 OAI21xp33_ASAP7_75t_R n_9325 (.A1(net19),
    .A2(n_8926_o_0),
    .B(n_9033_o_0),
    .Y(n_9325_o_0));
 AO22x1_ASAP7_75t_R n_9326 (.A1(n_9165_o_0),
    .A2(n_9324_o_0),
    .B1(n_9325_o_0),
    .B2(n_8942_o_0),
    .Y(n_9326_o_0));
 NAND2xp33_ASAP7_75t_R n_9327 (.A(n_9229_o_0),
    .B(n_9010_o_0),
    .Y(n_9327_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9328 (.A1(n_8926_o_0),
    .A2(n_9077_o_0),
    .B(n_9027_o_0),
    .C(n_9327_o_0),
    .Y(n_9328_o_0));
 AOI211xp5_ASAP7_75t_R n_9329 (.A1(n_8889_o_0),
    .A2(n_9326_o_0),
    .B(n_9328_o_0),
    .C(n_9024_o_0),
    .Y(n_9329_o_0));
 INVx1_ASAP7_75t_R n_933 (.A(n_847_o_0),
    .Y(n_933_o_0));
 AOI21xp33_ASAP7_75t_R n_9330 (.A1(n_9178_o_0),
    .A2(n_9323_o_0),
    .B(n_9329_o_0),
    .Y(n_9330_o_0));
 INVx1_ASAP7_75t_R n_9331 (.A(n_9324_o_0),
    .Y(n_9331_o_0));
 NAND3xp33_ASAP7_75t_R n_9332 (.A(n_8995_o_0),
    .B(n_9040_o_0),
    .C(n_8942_o_0),
    .Y(n_9332_o_0));
 OAI31xp33_ASAP7_75t_R n_9333 (.A1(n_9146_o_0),
    .A2(n_9331_o_0),
    .A3(n_8942_o_0),
    .B(n_9332_o_0),
    .Y(n_9333_o_0));
 NAND3xp33_ASAP7_75t_R n_9334 (.A(n_9001_o_0),
    .B(n_9024_o_0),
    .C(n_8942_o_0),
    .Y(n_9334_o_0));
 INVx1_ASAP7_75t_R n_9335 (.A(n_8959_o_0),
    .Y(n_9335_o_0));
 OAI221xp5_ASAP7_75t_R n_9336 (.A1(n_9334_o_0),
    .A2(n_8970_o_0),
    .B1(n_9046_o_0),
    .B2(n_9335_o_0),
    .C(net64),
    .Y(n_9336_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9337 (.A1(n_8968_o_0),
    .A2(n_9140_o_0),
    .B(n_9106_o_0),
    .C(n_9041_o_0),
    .Y(n_9337_o_0));
 OAI211xp5_ASAP7_75t_R n_9338 (.A1(net19),
    .A2(n_8926_o_0),
    .B(n_9024_o_0),
    .C(n_8942_o_0),
    .Y(n_9338_o_0));
 AOI211xp5_ASAP7_75t_R n_9339 (.A1(n_9315_o_0),
    .A2(n_9338_o_0),
    .B(n_8976_o_0),
    .C(n_9046_o_0),
    .Y(n_9339_o_0));
 NOR2xp33_ASAP7_75t_R n_934 (.A(n_836_o_0),
    .B(n_933_o_0),
    .Y(n_934_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9340 (.A1(n_8993_o_0),
    .A2(n_9337_o_0),
    .B(n_9339_o_0),
    .C(n_9010_o_0),
    .Y(n_9340_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9341 (.A1(n_8993_o_0),
    .A2(n_9333_o_0),
    .B(n_9336_o_0),
    .C(n_9340_o_0),
    .Y(n_9341_o_0));
 OAI22xp33_ASAP7_75t_R n_9342 (.A1(n_9330_o_0),
    .A2(n_8984_o_0),
    .B1(n_9008_o_0),
    .B2(n_9341_o_0),
    .Y(n_9342_o_0));
 NOR2xp33_ASAP7_75t_R n_9343 (.A(n_8926_o_0),
    .B(n_8960_o_0),
    .Y(n_9343_o_0));
 OAI21xp33_ASAP7_75t_R n_9344 (.A1(n_8963_o_0),
    .A2(n_9001_o_0),
    .B(n_9010_o_0),
    .Y(n_9344_o_0));
 AOI21xp33_ASAP7_75t_R n_9345 (.A1(n_9093_o_0),
    .A2(n_8946_o_0),
    .B(n_9344_o_0),
    .Y(n_9345_o_0));
 OA21x2_ASAP7_75t_R n_9346 (.A1(n_8998_o_0),
    .A2(n_9343_o_0),
    .B(n_9345_o_0),
    .Y(n_9346_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9347 (.A1(net19),
    .A2(n_8946_o_0),
    .B(n_8926_o_0),
    .C(n_8942_o_0),
    .Y(n_9347_o_0));
 INVx1_ASAP7_75t_R n_9348 (.A(n_9347_o_0),
    .Y(n_9348_o_0));
 AOI321xp33_ASAP7_75t_R n_9349 (.A1(n_8939_o_0),
    .A2(n_9054_o_0),
    .A3(n_8926_o_0),
    .B1(n_9093_o_0),
    .B2(n_9077_o_0),
    .C(n_9037_o_0),
    .Y(n_9349_o_0));
 NAND2xp5_ASAP7_75t_R n_935 (.A(n_847_o_0),
    .B(n_864_o_0),
    .Y(n_935_o_0));
 OA21x2_ASAP7_75t_R n_9350 (.A1(n_9348_o_0),
    .A2(n_8927_o_0),
    .B(n_9349_o_0),
    .Y(n_9350_o_0));
 AOI21xp33_ASAP7_75t_R n_9351 (.A1(n_8958_o_0),
    .A2(n_9033_o_0),
    .B(n_8968_o_0),
    .Y(n_9351_o_0));
 NOR2xp33_ASAP7_75t_R n_9352 (.A(n_8942_o_0),
    .B(n_8974_o_0),
    .Y(n_9352_o_0));
 AO21x1_ASAP7_75t_R n_9353 (.A1(n_9093_o_0),
    .A2(n_9054_o_0),
    .B(n_8949_o_0),
    .Y(n_9353_o_0));
 OAI321xp33_ASAP7_75t_R n_9354 (.A1(n_9010_o_0),
    .A2(n_9351_o_0),
    .A3(n_9352_o_0),
    .B1(n_9353_o_0),
    .B2(n_9344_o_0),
    .C(n_8993_o_0),
    .Y(n_9354_o_0));
 OAI31xp33_ASAP7_75t_R n_9355 (.A1(n_9046_o_0),
    .A2(n_9346_o_0),
    .A3(n_9350_o_0),
    .B(n_9354_o_0),
    .Y(n_9355_o_0));
 INVx1_ASAP7_75t_R n_9356 (.A(n_9035_o_0),
    .Y(n_9356_o_0));
 AOI31xp33_ASAP7_75t_R n_9357 (.A1(n_8939_o_0),
    .A2(n_9043_o_0),
    .A3(n_9040_o_0),
    .B(n_8993_o_0),
    .Y(n_9357_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9358 (.A1(n_8926_o_0),
    .A2(n_8915_o_0),
    .B(n_9356_o_0),
    .C(n_9357_o_0),
    .Y(n_9358_o_0));
 OA21x2_ASAP7_75t_R n_9359 (.A1(n_8978_o_0),
    .A2(n_9120_o_0),
    .B(n_9046_o_0),
    .Y(n_9359_o_0));
 OAI21xp33_ASAP7_75t_R n_936 (.A1(n_881_o_0),
    .A2(n_935_o_0),
    .B(n_877_o_0),
    .Y(n_936_o_0));
 OAI21xp33_ASAP7_75t_R n_9360 (.A1(n_9335_o_0),
    .A2(n_9060_o_0),
    .B(n_9359_o_0),
    .Y(n_9360_o_0));
 AOI21xp33_ASAP7_75t_R n_9361 (.A1(n_9358_o_0),
    .A2(n_9360_o_0),
    .B(n_9010_o_0),
    .Y(n_9361_o_0));
 INVx1_ASAP7_75t_R n_9362 (.A(n_9149_o_0),
    .Y(n_9362_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9363 (.A1(n_8915_o_0),
    .A2(n_8926_o_0),
    .B(net19),
    .C(n_8939_o_0),
    .Y(n_9363_o_0));
 OAI31xp33_ASAP7_75t_R n_9364 (.A1(n_8939_o_0),
    .A2(n_9133_o_0),
    .A3(n_8926_o_0),
    .B(n_9363_o_0),
    .Y(n_9364_o_0));
 AOI21xp33_ASAP7_75t_R n_9365 (.A1(n_9024_o_0),
    .A2(n_9364_o_0),
    .B(n_8889_o_0),
    .Y(n_9365_o_0));
 OA21x2_ASAP7_75t_R n_9366 (.A1(n_9362_o_0),
    .A2(n_9196_o_0),
    .B(n_9365_o_0),
    .Y(n_9366_o_0));
 OAI21xp33_ASAP7_75t_R n_9367 (.A1(n_9361_o_0),
    .A2(n_9366_o_0),
    .B(n_8983_o_0),
    .Y(n_9367_o_0));
 OAI211xp5_ASAP7_75t_R n_9368 (.A1(n_9008_o_0),
    .A2(n_9355_o_0),
    .B(n_9367_o_0),
    .C(n_8872_o_0),
    .Y(n_9368_o_0));
 OAI21xp33_ASAP7_75t_R n_9369 (.A1(n_9105_o_0),
    .A2(n_9342_o_0),
    .B(n_9368_o_0),
    .Y(n_9369_o_0));
 AOI21xp33_ASAP7_75t_R n_937 (.A1(n_881_o_0),
    .A2(n_889_o_0),
    .B(n_877_o_0),
    .Y(n_937_o_0));
 NOR3xp33_ASAP7_75t_R n_9370 (.A(n_9006_o_0),
    .B(n_8970_o_0),
    .C(n_8939_o_0),
    .Y(n_9370_o_0));
 AOI31xp33_ASAP7_75t_R n_9371 (.A1(n_8942_o_0),
    .A2(n_8979_o_0),
    .A3(n_9072_o_0),
    .B(n_9370_o_0),
    .Y(n_9371_o_0));
 AO21x1_ASAP7_75t_R n_9372 (.A1(n_8928_o_0),
    .A2(n_9347_o_0),
    .B(n_9137_o_0),
    .Y(n_9372_o_0));
 AOI21xp33_ASAP7_75t_R n_9373 (.A1(n_8972_o_0),
    .A2(n_9372_o_0),
    .B(n_9046_o_0),
    .Y(n_9373_o_0));
 AOI22xp33_ASAP7_75t_R n_9374 (.A1(n_9093_o_0),
    .A2(n_9077_o_0),
    .B1(n_8939_o_0),
    .B2(n_9039_o_0),
    .Y(n_9374_o_0));
 OAI21xp33_ASAP7_75t_R n_9375 (.A1(n_9011_o_0),
    .A2(n_9056_o_0),
    .B(n_9374_o_0),
    .Y(n_9375_o_0));
 AOI21xp33_ASAP7_75t_R n_9376 (.A1(n_9106_o_0),
    .A2(n_9237_o_0),
    .B(n_9037_o_0),
    .Y(n_9376_o_0));
 AOI211xp5_ASAP7_75t_R n_9377 (.A1(n_9375_o_0),
    .A2(n_9037_o_0),
    .B(n_8992_o_0),
    .C(n_9376_o_0),
    .Y(n_9377_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9378 (.A1(net64),
    .A2(n_9371_o_0),
    .B(n_9373_o_0),
    .C(n_9377_o_0),
    .Y(n_9378_o_0));
 NAND2xp33_ASAP7_75t_R n_9379 (.A(n_9324_o_0),
    .B(n_9004_o_0),
    .Y(n_9379_o_0));
 NOR2xp33_ASAP7_75t_R n_938 (.A(n_881_o_0),
    .B(n_913_o_0),
    .Y(n_938_o_0));
 OAI31xp33_ASAP7_75t_R n_9380 (.A1(n_8968_o_0),
    .A2(n_9140_o_0),
    .A3(n_9131_o_0),
    .B(n_9379_o_0),
    .Y(n_9380_o_0));
 OAI21xp33_ASAP7_75t_R n_9381 (.A1(n_8915_o_0),
    .A2(n_8942_o_0),
    .B(n_9010_o_0),
    .Y(n_9381_o_0));
 AOI21xp33_ASAP7_75t_R n_9382 (.A1(n_8974_o_0),
    .A2(n_8947_o_0),
    .B(n_9063_o_0),
    .Y(n_9382_o_0));
 OAI21xp33_ASAP7_75t_R n_9383 (.A1(n_9381_o_0),
    .A2(n_9382_o_0),
    .B(n_9046_o_0),
    .Y(n_9383_o_0));
 AOI21xp33_ASAP7_75t_R n_9384 (.A1(n_8889_o_0),
    .A2(n_9380_o_0),
    .B(n_9383_o_0),
    .Y(n_9384_o_0));
 OAI22xp33_ASAP7_75t_R n_9385 (.A1(n_9335_o_0),
    .A2(n_9005_o_0),
    .B1(n_8963_o_0),
    .B2(n_9056_o_0),
    .Y(n_9385_o_0));
 OAI31xp33_ASAP7_75t_R n_9386 (.A1(n_9037_o_0),
    .A2(n_9282_o_0),
    .A3(n_9214_o_0),
    .B(n_8992_o_0),
    .Y(n_9386_o_0));
 AOI21xp33_ASAP7_75t_R n_9387 (.A1(n_9010_o_0),
    .A2(n_9385_o_0),
    .B(n_9386_o_0),
    .Y(n_9387_o_0));
 OAI21xp33_ASAP7_75t_R n_9388 (.A1(n_9384_o_0),
    .A2(n_9387_o_0),
    .B(n_8983_o_0),
    .Y(n_9388_o_0));
 OAI21xp33_ASAP7_75t_R n_9389 (.A1(n_8983_o_0),
    .A2(n_9378_o_0),
    .B(n_9388_o_0),
    .Y(n_9389_o_0));
 INVx1_ASAP7_75t_R n_939 (.A(n_938_o_0),
    .Y(n_939_o_0));
 AOI31xp33_ASAP7_75t_R n_9390 (.A1(net19),
    .A2(n_8947_o_0),
    .A3(n_8968_o_0),
    .B(n_9111_o_0),
    .Y(n_9390_o_0));
 OA21x2_ASAP7_75t_R n_9391 (.A1(n_8968_o_0),
    .A2(n_9078_o_0),
    .B(n_9038_o_0),
    .Y(n_9391_o_0));
 AOI211xp5_ASAP7_75t_R n_9392 (.A1(n_9390_o_0),
    .A2(n_9238_o_0),
    .B(n_8992_o_0),
    .C(n_9391_o_0),
    .Y(n_9392_o_0));
 OAI21xp33_ASAP7_75t_R n_9393 (.A1(n_8947_o_0),
    .A2(n_8960_o_0),
    .B(n_8942_o_0),
    .Y(n_9393_o_0));
 OAI22xp33_ASAP7_75t_R n_9394 (.A1(n_9073_o_0),
    .A2(n_9393_o_0),
    .B1(n_9011_o_0),
    .B2(n_9034_o_0),
    .Y(n_9394_o_0));
 AOI321xp33_ASAP7_75t_R n_9395 (.A1(n_8963_o_0),
    .A2(n_9072_o_0),
    .A3(n_9001_o_0),
    .B1(n_8942_o_0),
    .B2(n_9124_o_0),
    .C(n_9010_o_0),
    .Y(n_9395_o_0));
 AOI21xp33_ASAP7_75t_R n_9396 (.A1(n_9037_o_0),
    .A2(n_9394_o_0),
    .B(n_9395_o_0),
    .Y(n_9396_o_0));
 OAI21xp33_ASAP7_75t_R n_9397 (.A1(n_9046_o_0),
    .A2(n_9396_o_0),
    .B(n_8983_o_0),
    .Y(n_9397_o_0));
 OAI21xp33_ASAP7_75t_R n_9398 (.A1(n_8942_o_0),
    .A2(n_9029_o_0),
    .B(n_9010_o_0),
    .Y(n_9398_o_0));
 AOI211xp5_ASAP7_75t_R n_9399 (.A1(n_8889_o_0),
    .A2(n_8974_o_0),
    .B(n_8926_o_0),
    .C(n_8968_o_0),
    .Y(n_9399_o_0));
 AOI21xp33_ASAP7_75t_R n_940 (.A1(n_937_o_0),
    .A2(n_939_o_0),
    .B(net14),
    .Y(n_940_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9400 (.A1(n_8968_o_0),
    .A2(n_9002_o_0),
    .B(n_9037_o_0),
    .C(n_9094_o_0),
    .D(n_9399_o_0),
    .Y(n_9400_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9401 (.A1(n_8947_o_0),
    .A2(n_9054_o_0),
    .B(n_9400_o_0),
    .C(n_9046_o_0),
    .Y(n_9401_o_0));
 OAI21xp33_ASAP7_75t_R n_9402 (.A1(n_9351_o_0),
    .A2(n_9398_o_0),
    .B(n_9401_o_0),
    .Y(n_9402_o_0));
 AOI21xp33_ASAP7_75t_R n_9403 (.A1(n_8947_o_0),
    .A2(n_9089_o_0),
    .B(n_8949_o_0),
    .Y(n_9403_o_0));
 OAI21xp33_ASAP7_75t_R n_9404 (.A1(n_9049_o_0),
    .A2(n_9393_o_0),
    .B(n_9403_o_0),
    .Y(n_9404_o_0));
 AOI21xp33_ASAP7_75t_R n_9405 (.A1(n_9165_o_0),
    .A2(n_9153_o_0),
    .B(n_8889_o_0),
    .Y(n_9405_o_0));
 OAI31xp33_ASAP7_75t_R n_9406 (.A1(n_8939_o_0),
    .A2(n_9005_o_0),
    .A3(n_9131_o_0),
    .B(n_9405_o_0),
    .Y(n_9406_o_0));
 OAI211xp5_ASAP7_75t_R n_9407 (.A1(n_9404_o_0),
    .A2(n_9010_o_0),
    .B(n_8993_o_0),
    .C(n_9406_o_0),
    .Y(n_9407_o_0));
 AOI31xp33_ASAP7_75t_R n_9408 (.A1(n_8880_o_0),
    .A2(n_9402_o_0),
    .A3(n_9407_o_0),
    .B(n_8873_o_0),
    .Y(n_9408_o_0));
 OAI21xp33_ASAP7_75t_R n_9409 (.A1(n_9392_o_0),
    .A2(n_9397_o_0),
    .B(n_9408_o_0),
    .Y(n_9409_o_0));
 NAND2xp33_ASAP7_75t_R n_941 (.A(n_881_o_0),
    .B(n_935_o_0),
    .Y(n_941_o_0));
 OAI21xp33_ASAP7_75t_R n_9410 (.A1(n_9105_o_0),
    .A2(n_9389_o_0),
    .B(n_9409_o_0),
    .Y(n_9410_o_0));
 NAND2xp33_ASAP7_75t_R n_9411 (.A(n_4959_o_0),
    .B(n_4823_o_0),
    .Y(n_9411_o_0));
 OAI21xp33_ASAP7_75t_R n_9412 (.A1(n_4823_o_0),
    .A2(n_4959_o_0),
    .B(n_9411_o_0),
    .Y(n_9412_o_0));
 NOR2xp33_ASAP7_75t_R n_9413 (.A(_01112_),
    .B(n_9412_o_0),
    .Y(n_9413_o_0));
 NOR2xp33_ASAP7_75t_R n_9414 (.A(_00721_),
    .B(net),
    .Y(n_9414_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9415 (.A1(n_9412_o_0),
    .A2(_01112_),
    .B(n_9413_o_0),
    .C(net),
    .D(n_9414_o_0),
    .Y(n_9415_o_0));
 HAxp5_ASAP7_75t_R n_9416 (.A(n_1422_o_0),
    .B(n_9415_o_0),
    .CON(n_9416_o_0),
    .SN(n_9416_o_1));
 INVx1_ASAP7_75t_R n_9417 (.A(n_9416_o_1),
    .Y(n_9417_o_0));
 XNOR2xp5_ASAP7_75t_R n_9418 (.A(_01113_),
    .B(n_4804_o_0),
    .Y(n_9418_o_0));
 NOR2xp33_ASAP7_75t_R n_9419 (.A(n_4812_o_0),
    .B(n_9418_o_0),
    .Y(n_9419_o_0));
 OAI21xp33_ASAP7_75t_R n_942 (.A1(n_881_o_0),
    .A2(n_935_o_0),
    .B(n_878_o_0),
    .Y(n_942_o_0));
 NOR2xp33_ASAP7_75t_R n_9420 (.A(_00720_),
    .B(net),
    .Y(n_9420_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9421 (.A1(n_4812_o_0),
    .A2(n_9418_o_0),
    .B(n_9419_o_0),
    .C(net),
    .D(n_9420_o_0),
    .Y(n_9421_o_0));
 XNOR2xp5_ASAP7_75t_R n_9422 (.A(_00970_),
    .B(n_9421_o_0),
    .Y(n_9422_o_0));
 INVx1_ASAP7_75t_R n_9423 (.A(_00966_),
    .Y(n_9423_o_0));
 XNOR2xp5_ASAP7_75t_R n_9424 (.A(_01022_),
    .B(_01030_),
    .Y(n_9424_o_0));
 NAND2xp33_ASAP7_75t_R n_9425 (.A(_01109_),
    .B(n_9424_o_0),
    .Y(n_9425_o_0));
 OAI21xp33_ASAP7_75t_R n_9426 (.A1(_01109_),
    .A2(n_9424_o_0),
    .B(n_9425_o_0),
    .Y(n_9426_o_0));
 OAI211xp5_ASAP7_75t_R n_9427 (.A1(_01109_),
    .A2(n_9424_o_0),
    .B(n_9425_o_0),
    .C(n_7158_o_0),
    .Y(n_9427_o_0));
 INVx1_ASAP7_75t_R n_9428 (.A(n_9427_o_0),
    .Y(n_9428_o_0));
 NOR2xp33_ASAP7_75t_R n_9429 (.A(_00608_),
    .B(_00858_),
    .Y(n_9429_o_0));
 INVx1_ASAP7_75t_R n_943 (.A(n_942_o_0),
    .Y(n_943_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9430 (.A1(n_7153_o_0),
    .A2(n_9426_o_0),
    .B(n_9428_o_0),
    .C(net39),
    .D(n_9429_o_0),
    .Y(n_9430_o_0));
 NOR2xp33_ASAP7_75t_R n_9431 (.A(_01109_),
    .B(n_9424_o_0),
    .Y(n_9431_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9432 (.A1(_01109_),
    .A2(n_9424_o_0),
    .B(n_9431_o_0),
    .C(n_7153_o_0),
    .Y(n_9432_o_0));
 INVx1_ASAP7_75t_R n_9433 (.A(n_9429_o_0),
    .Y(n_9433_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9434 (.A1(n_9427_o_0),
    .A2(n_9432_o_0),
    .B(n_3021_o_0),
    .C(n_9433_o_0),
    .D(n_9423_o_0),
    .Y(n_9434_o_0));
 AOI21x1_ASAP7_75t_R n_9435 (.A1(n_9423_o_0),
    .A2(n_9430_o_0),
    .B(n_9434_o_0),
    .Y(n_9435_o_0));
 NAND2xp33_ASAP7_75t_R n_9436 (.A(_01107_),
    .B(_01114_),
    .Y(n_9436_o_0));
 OAI21xp33_ASAP7_75t_R n_9437 (.A1(_01107_),
    .A2(_01114_),
    .B(n_9436_o_0),
    .Y(n_9437_o_0));
 XNOR2xp5_ASAP7_75t_R n_9438 (.A(_01028_),
    .B(_01075_),
    .Y(n_9438_o_0));
 NAND2xp33_ASAP7_75t_R n_9439 (.A(n_4922_o_0),
    .B(n_9438_o_0),
    .Y(n_9439_o_0));
 NAND2xp33_ASAP7_75t_R n_944 (.A(n_847_o_0),
    .B(n_836_o_0),
    .Y(n_944_o_0));
 OAI21xp33_ASAP7_75t_R n_9440 (.A1(n_9438_o_0),
    .A2(n_4922_o_0),
    .B(n_9439_o_0),
    .Y(n_9440_o_0));
 NOR2xp33_ASAP7_75t_R n_9441 (.A(n_4922_o_0),
    .B(n_9438_o_0),
    .Y(n_9441_o_0));
 AOI211xp5_ASAP7_75t_R n_9442 (.A1(n_9438_o_0),
    .A2(n_4922_o_0),
    .B(n_9441_o_0),
    .C(n_9437_o_0),
    .Y(n_9442_o_0));
 NOR2xp33_ASAP7_75t_R n_9443 (.A(_00606_),
    .B(_00858_),
    .Y(n_9443_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9444 (.A1(n_9437_o_0),
    .A2(n_9440_o_0),
    .B(n_9442_o_0),
    .C(net77),
    .D(n_9443_o_0),
    .Y(n_9444_o_0));
 NOR2xp33_ASAP7_75t_R n_9445 (.A(_01107_),
    .B(_01114_),
    .Y(n_9445_o_0));
 AOI21xp33_ASAP7_75t_R n_9446 (.A1(_01107_),
    .A2(_01114_),
    .B(n_9445_o_0),
    .Y(n_9446_o_0));
 OAI211xp5_ASAP7_75t_R n_9447 (.A1(n_9438_o_0),
    .A2(n_4922_o_0),
    .B(n_9439_o_0),
    .C(n_9446_o_0),
    .Y(n_9447_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9448 (.A1(n_9438_o_0),
    .A2(n_4922_o_0),
    .B(n_9441_o_0),
    .C(n_9437_o_0),
    .Y(n_9448_o_0));
 INVx1_ASAP7_75t_R n_9449 (.A(n_9443_o_0),
    .Y(n_9449_o_0));
 INVx1_ASAP7_75t_R n_945 (.A(n_944_o_0),
    .Y(n_945_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9450 (.A1(n_9447_o_0),
    .A2(n_9448_o_0),
    .B(net3),
    .C(n_9449_o_0),
    .D(_00964_),
    .Y(n_9450_o_0));
 AOI21x1_ASAP7_75t_R n_9451 (.A1(_00964_),
    .A2(n_9444_o_0),
    .B(n_9450_o_0),
    .Y(n_9451_o_0));
 INVx1_ASAP7_75t_R n_9452 (.A(n_9451_o_0),
    .Y(n_9452_o_0));
 NAND2xp33_ASAP7_75t_R n_9453 (.A(n_9435_o_0),
    .B(n_9452_o_0),
    .Y(n_9453_o_0));
 NOR2xp33_ASAP7_75t_R n_9454 (.A(_00723_),
    .B(_00858_),
    .Y(n_9454_o_0));
 XNOR2xp5_ASAP7_75t_R n_9455 (.A(_01023_),
    .B(_01031_),
    .Y(n_9455_o_0));
 XNOR2xp5_ASAP7_75t_R n_9456 (.A(_01109_),
    .B(_01114_),
    .Y(n_9456_o_0));
 NAND2xp33_ASAP7_75t_R n_9457 (.A(n_9455_o_0),
    .B(n_9456_o_0),
    .Y(n_9457_o_0));
 OAI21xp33_ASAP7_75t_R n_9458 (.A1(n_9455_o_0),
    .A2(n_9456_o_0),
    .B(n_9457_o_0),
    .Y(n_9458_o_0));
 NAND2xp33_ASAP7_75t_R n_9459 (.A(_01110_),
    .B(n_7143_o_0),
    .Y(n_9459_o_0));
 OAI21xp33_ASAP7_75t_R n_946 (.A1(n_878_o_0),
    .A2(n_945_o_0),
    .B(n_891_o_0),
    .Y(n_946_o_0));
 OAI21xp33_ASAP7_75t_R n_9460 (.A1(_01110_),
    .A2(n_7143_o_0),
    .B(n_9459_o_0),
    .Y(n_9460_o_0));
 NAND2xp33_ASAP7_75t_R n_9461 (.A(n_9458_o_0),
    .B(n_9460_o_0),
    .Y(n_9461_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9462 (.A1(n_9458_o_0),
    .A2(n_9460_o_0),
    .B(n_9461_o_0),
    .C(n_3021_o_0),
    .Y(n_9462_o_0));
 INVx1_ASAP7_75t_R n_9463 (.A(_00967_),
    .Y(n_9463_o_0));
 OAI21xp33_ASAP7_75t_R n_9464 (.A1(n_9454_o_0),
    .A2(n_9462_o_0),
    .B(n_9463_o_0),
    .Y(n_9464_o_0));
 OAI31xp33_ASAP7_75t_R n_9465 (.A1(n_9454_o_0),
    .A2(n_9462_o_0),
    .A3(n_9463_o_0),
    .B(n_9464_o_0),
    .Y(n_9465_o_0));
 NAND2xp33_ASAP7_75t_R n_9466 (.A(n_7152_o_0),
    .B(n_9446_o_0),
    .Y(n_9466_o_0));
 OAI21xp33_ASAP7_75t_R n_9467 (.A1(n_7152_o_0),
    .A2(n_9446_o_0),
    .B(n_9466_o_0),
    .Y(n_9467_o_0));
 OAI211xp5_ASAP7_75t_R n_9468 (.A1(_01021_),
    .A2(_01029_),
    .B(n_4860_o_0),
    .C(n_4901_o_0),
    .Y(n_9468_o_0));
 OAI21xp33_ASAP7_75t_R n_9469 (.A1(n_4901_o_0),
    .A2(n_4862_o_0),
    .B(n_9468_o_0),
    .Y(n_9469_o_0));
 AOI21xp33_ASAP7_75t_R n_947 (.A1(n_941_o_0),
    .A2(n_943_o_0),
    .B(n_946_o_0),
    .Y(n_947_o_0));
 NOR2xp33_ASAP7_75t_R n_9470 (.A(n_9437_o_0),
    .B(n_7156_o_0),
    .Y(n_9470_o_0));
 NOR2xp33_ASAP7_75t_R n_9471 (.A(n_7152_o_0),
    .B(n_9446_o_0),
    .Y(n_9471_o_0));
 OAI21xp33_ASAP7_75t_R n_9472 (.A1(n_9470_o_0),
    .A2(n_9471_o_0),
    .B(n_9469_o_0),
    .Y(n_9472_o_0));
 OAI211xp5_ASAP7_75t_R n_9473 (.A1(n_9467_o_0),
    .A2(n_9469_o_0),
    .B(n_9472_o_0),
    .C(net39),
    .Y(n_9473_o_0));
 NAND2xp33_ASAP7_75t_R n_9474 (.A(_00605_),
    .B(n_3021_o_0),
    .Y(n_9474_o_0));
 INVx1_ASAP7_75t_R n_9475 (.A(_00965_),
    .Y(n_9475_o_0));
 INVx1_ASAP7_75t_R n_9476 (.A(_00605_),
    .Y(n_9476_o_0));
 INVx1_ASAP7_75t_R n_9477 (.A(n_9445_o_0),
    .Y(n_9477_o_0));
 XNOR2xp5_ASAP7_75t_R n_9478 (.A(n_4901_o_0),
    .B(n_4861_o_0),
    .Y(n_9478_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9479 (.A1(n_9477_o_0),
    .A2(n_9436_o_0),
    .B(n_7152_o_0),
    .C(n_9466_o_0),
    .D(n_9478_o_0),
    .Y(n_9479_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_948 (.A1(n_934_o_0),
    .A2(n_936_o_0),
    .B(n_940_o_0),
    .C(n_947_o_0),
    .Y(n_948_o_0));
 OAI31xp33_ASAP7_75t_R n_9480 (.A1(n_9470_o_0),
    .A2(n_9469_o_0),
    .A3(n_9471_o_0),
    .B(net39),
    .Y(n_9480_o_0));
 OAI221xp5_ASAP7_75t_R n_9481 (.A1(net39),
    .A2(n_9476_o_0),
    .B1(n_9479_o_0),
    .B2(n_9480_o_0),
    .C(n_9475_o_0),
    .Y(n_9481_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9482 (.A1(n_9473_o_0),
    .A2(n_9474_o_0),
    .B(n_9475_o_0),
    .C(n_9481_o_0),
    .Y(n_9482_o_0));
 NOR2xp33_ASAP7_75t_R n_9483 (.A(n_9482_o_0),
    .B(n_9451_o_0),
    .Y(n_9483_o_0));
 INVx1_ASAP7_75t_R n_9484 (.A(_00723_),
    .Y(n_9484_o_0));
 AOI21xp33_ASAP7_75t_R n_9485 (.A1(n_9484_o_0),
    .A2(net3),
    .B(n_9462_o_0),
    .Y(n_9485_o_0));
 XNOR2xp5_ASAP7_75t_R n_9486 (.A(_01110_),
    .B(n_7137_o_0),
    .Y(n_9486_o_0));
 XNOR2xp5_ASAP7_75t_R n_9487 (.A(n_9486_o_0),
    .B(n_9458_o_0),
    .Y(n_9487_o_0));
 INVx1_ASAP7_75t_R n_9488 (.A(n_9454_o_0),
    .Y(n_9488_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9489 (.A1(net1),
    .A2(n_9487_o_0),
    .B(n_9488_o_0),
    .C(_00967_),
    .Y(n_9489_o_0));
 NOR2xp33_ASAP7_75t_R n_949 (.A(net32),
    .B(n_913_o_0),
    .Y(n_949_o_0));
 AOI21xp5_ASAP7_75t_R n_9490 (.A1(_00967_),
    .A2(n_9485_o_0),
    .B(n_9489_o_0),
    .Y(n_9490_o_0));
 OAI21xp33_ASAP7_75t_R n_9491 (.A1(n_9435_o_0),
    .A2(net22),
    .B(n_9490_o_0),
    .Y(n_9491_o_0));
 NAND2xp33_ASAP7_75t_R n_9492 (.A(n_9435_o_0),
    .B(n_9483_o_0),
    .Y(n_9492_o_0));
 INVx1_ASAP7_75t_R n_9493 (.A(n_9492_o_0),
    .Y(n_9493_o_0));
 XNOR2xp5_ASAP7_75t_R n_9494 (.A(_01111_),
    .B(n_7208_o_0),
    .Y(n_9494_o_0));
 XNOR2xp5_ASAP7_75t_R n_9495 (.A(_01110_),
    .B(_01114_),
    .Y(n_9495_o_0));
 XNOR2xp5_ASAP7_75t_R n_9496 (.A(n_4802_o_0),
    .B(n_9495_o_0),
    .Y(n_9496_o_0));
 XOR2xp5_ASAP7_75t_R n_9497 (.A(n_9494_o_0),
    .B(n_9496_o_0),
    .Y(n_9497_o_0));
 NOR2xp33_ASAP7_75t_R n_9498 (.A(_00722_),
    .B(net39),
    .Y(n_9498_o_0));
 AOI21xp33_ASAP7_75t_R n_9499 (.A1(net),
    .A2(n_9497_o_0),
    .B(n_9498_o_0),
    .Y(n_9499_o_0));
 INVx1_ASAP7_75t_R n_950 (.A(n_949_o_0),
    .Y(n_950_o_0));
 NOR2xp33_ASAP7_75t_R n_9500 (.A(n_1359_o_0),
    .B(n_9499_o_0),
    .Y(n_9500_o_0));
 AOI21xp33_ASAP7_75t_R n_9501 (.A1(n_1359_o_0),
    .A2(n_9499_o_0),
    .B(n_9500_o_0),
    .Y(n_9501_o_0));
 OAI21xp33_ASAP7_75t_R n_9502 (.A1(n_9491_o_0),
    .A2(n_9493_o_0),
    .B(n_9501_o_0),
    .Y(n_9502_o_0));
 AOI21xp33_ASAP7_75t_R n_9503 (.A1(n_9453_o_0),
    .A2(n_9465_o_0),
    .B(n_9502_o_0),
    .Y(n_9503_o_0));
 AOI21xp33_ASAP7_75t_R n_9504 (.A1(n_9435_o_0),
    .A2(n_9483_o_0),
    .B(n_9490_o_0),
    .Y(n_9504_o_0));
 NOR2xp33_ASAP7_75t_R n_9505 (.A(n_9451_o_0),
    .B(n_9435_o_0),
    .Y(n_9505_o_0));
 INVx1_ASAP7_75t_R n_9506 (.A(n_9505_o_0),
    .Y(n_9506_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9507 (.A1(net1),
    .A2(n_9487_o_0),
    .B(n_9488_o_0),
    .C(n_9463_o_0),
    .Y(n_9507_o_0));
 AOI21x1_ASAP7_75t_R n_9508 (.A1(n_9463_o_0),
    .A2(n_9485_o_0),
    .B(n_9507_o_0),
    .Y(n_9508_o_0));
 OAI21xp33_ASAP7_75t_R n_9509 (.A1(net53),
    .A2(n_9452_o_0),
    .B(n_9435_o_0),
    .Y(n_9509_o_0));
 NAND3xp33_ASAP7_75t_R n_951 (.A(n_950_o_0),
    .B(n_944_o_0),
    .C(n_878_o_0),
    .Y(n_951_o_0));
 INVx1_ASAP7_75t_R n_9510 (.A(n_9509_o_0),
    .Y(n_9510_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9511 (.A1(_00964_),
    .A2(n_9444_o_0),
    .B(n_9450_o_0),
    .C(n_9482_o_0),
    .Y(n_9511_o_0));
 INVx1_ASAP7_75t_R n_9512 (.A(n_9473_o_0),
    .Y(n_9512_o_0));
 INVx1_ASAP7_75t_R n_9513 (.A(n_9474_o_0),
    .Y(n_9513_o_0));
 INVx1_ASAP7_75t_R n_9514 (.A(n_9468_o_0),
    .Y(n_9514_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9515 (.A1(n_4861_o_0),
    .A2(_01108_),
    .B(n_9514_o_0),
    .C(net),
    .Y(n_9515_o_0));
 OAI21xp33_ASAP7_75t_R n_9516 (.A1(n_9470_o_0),
    .A2(n_9471_o_0),
    .B(net),
    .Y(n_9516_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9517 (.A1(n_9467_o_0),
    .A2(n_9515_o_0),
    .B(n_9516_o_0),
    .C(n_9479_o_0),
    .Y(n_9517_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9518 (.A1(net2),
    .A2(_00605_),
    .B(n_9517_o_0),
    .C(_00965_),
    .Y(n_9518_o_0));
 OAI311xp33_ASAP7_75t_R n_9519 (.A1(_00965_),
    .A2(n_9512_o_0),
    .A3(n_9513_o_0),
    .B1(n_9451_o_0),
    .C1(n_9518_o_0),
    .Y(n_9519_o_0));
 NOR2xp33_ASAP7_75t_R n_952 (.A(n_864_o_0),
    .B(n_836_o_0),
    .Y(n_952_o_0));
 AOI21xp33_ASAP7_75t_R n_9520 (.A1(n_9519_o_0),
    .A2(n_9511_o_0),
    .B(n_9435_o_0),
    .Y(n_9520_o_0));
 AOI211xp5_ASAP7_75t_R n_9521 (.A1(n_9497_o_0),
    .A2(net),
    .B(n_1359_o_0),
    .C(n_9498_o_0),
    .Y(n_9521_o_0));
 NOR2xp33_ASAP7_75t_R n_9522 (.A(_00968_),
    .B(n_9499_o_0),
    .Y(n_9522_o_0));
 NOR2xp67_ASAP7_75t_R n_9523 (.A(n_9521_o_0),
    .B(n_9522_o_0),
    .Y(n_9523_o_0));
 OAI31xp33_ASAP7_75t_R n_9524 (.A1(n_9508_o_0),
    .A2(n_9510_o_0),
    .A3(net85),
    .B(n_9523_o_0),
    .Y(n_9524_o_0));
 AOI21xp33_ASAP7_75t_R n_9525 (.A1(n_9504_o_0),
    .A2(n_9506_o_0),
    .B(n_9524_o_0),
    .Y(n_9525_o_0));
 INVx1_ASAP7_75t_R n_9526 (.A(n_9523_o_0),
    .Y(n_9526_o_0));
 NAND2xp33_ASAP7_75t_R n_9527 (.A(n_9482_o_0),
    .B(n_9452_o_0),
    .Y(n_9527_o_0));
 INVx1_ASAP7_75t_R n_9528 (.A(n_9527_o_0),
    .Y(n_9528_o_0));
 NOR2xp33_ASAP7_75t_R n_9529 (.A(n_9435_o_0),
    .B(n_9452_o_0),
    .Y(n_9529_o_0));
 INVx1_ASAP7_75t_R n_953 (.A(n_952_o_0),
    .Y(n_953_o_0));
 NOR3xp33_ASAP7_75t_R n_9530 (.A(n_9528_o_0),
    .B(n_9529_o_0),
    .C(n_9490_o_0),
    .Y(n_9530_o_0));
 AO21x1_ASAP7_75t_R n_9531 (.A1(n_9430_o_0),
    .A2(n_9423_o_0),
    .B(n_9434_o_0),
    .Y(n_9531_o_0));
 NAND2xp33_ASAP7_75t_R n_9532 (.A(n_9451_o_0),
    .B(n_9531_o_0),
    .Y(n_9532_o_0));
 AOI21xp33_ASAP7_75t_R n_9533 (.A1(n_9527_o_0),
    .A2(n_9532_o_0),
    .B(n_9465_o_0),
    .Y(n_9533_o_0));
 NAND3xp33_ASAP7_75t_R n_9534 (.A(n_9452_o_0),
    .B(net26),
    .C(n_9435_o_0),
    .Y(n_9534_o_0));
 INVx1_ASAP7_75t_R n_9535 (.A(n_9534_o_0),
    .Y(n_9535_o_0));
 NAND2xp33_ASAP7_75t_R n_9536 (.A(n_9427_o_0),
    .B(n_9432_o_0),
    .Y(n_9536_o_0));
 AOI211xp5_ASAP7_75t_R n_9537 (.A1(n_9536_o_0),
    .A2(net),
    .B(_00966_),
    .C(n_9429_o_0),
    .Y(n_9537_o_0));
 OAI211xp5_ASAP7_75t_R n_9538 (.A1(n_9537_o_0),
    .A2(n_9434_o_0),
    .B(net53),
    .C(n_9451_o_0),
    .Y(n_9538_o_0));
 INVx1_ASAP7_75t_R n_9539 (.A(n_9538_o_0),
    .Y(n_9539_o_0));
 INVx1_ASAP7_75t_R n_954 (.A(n_936_o_0),
    .Y(n_954_o_0));
 OAI221xp5_ASAP7_75t_R n_9540 (.A1(n_9452_o_0),
    .A2(net26),
    .B1(n_9435_o_0),
    .B2(net89),
    .C(n_9465_o_0),
    .Y(n_9540_o_0));
 OAI31xp33_ASAP7_75t_R n_9541 (.A1(n_9508_o_0),
    .A2(n_9535_o_0),
    .A3(n_9539_o_0),
    .B(n_9540_o_0),
    .Y(n_9541_o_0));
 XNOR2xp5_ASAP7_75t_R n_9542 (.A(n_1359_o_0),
    .B(n_9499_o_0),
    .Y(n_9542_o_0));
 NAND2xp33_ASAP7_75t_R n_9543 (.A(_00970_),
    .B(n_9421_o_0),
    .Y(n_9543_o_0));
 OAI21xp33_ASAP7_75t_R n_9544 (.A1(_00970_),
    .A2(n_9421_o_0),
    .B(n_9543_o_0),
    .Y(n_9544_o_0));
 OAI321xp33_ASAP7_75t_R n_9545 (.A1(n_9526_o_0),
    .A2(n_9530_o_0),
    .A3(n_9533_o_0),
    .B1(n_9541_o_0),
    .B2(n_9542_o_0),
    .C(n_9544_o_0),
    .Y(n_9545_o_0));
 OAI31xp33_ASAP7_75t_R n_9546 (.A1(n_9422_o_0),
    .A2(n_9503_o_0),
    .A3(n_9525_o_0),
    .B(n_9545_o_0),
    .Y(n_9546_o_0));
 XOR2xp5_ASAP7_75t_R n_9547 (.A(_01113_),
    .B(_01114_),
    .Y(n_9547_o_0));
 XNOR2xp5_ASAP7_75t_R n_9548 (.A(_01074_),
    .B(n_9547_o_0),
    .Y(n_9548_o_0));
 NOR2xp33_ASAP7_75t_R n_9549 (.A(n_4879_o_0),
    .B(n_9548_o_0),
    .Y(n_9549_o_0));
 AOI21xp33_ASAP7_75t_R n_955 (.A1(n_953_o_0),
    .A2(n_954_o_0),
    .B(net14),
    .Y(n_955_o_0));
 NOR2xp33_ASAP7_75t_R n_9550 (.A(_00719_),
    .B(net),
    .Y(n_9550_o_0));
 A2O1A1O1Ixp25_ASAP7_75t_R n_9551 (.A1(n_4879_o_0),
    .A2(n_9548_o_0),
    .B(n_9549_o_0),
    .C(net),
    .D(n_9550_o_0),
    .Y(n_9551_o_0));
 NAND2xp33_ASAP7_75t_R n_9552 (.A(_00971_),
    .B(n_9551_o_0),
    .Y(n_9552_o_0));
 OAI21xp33_ASAP7_75t_R n_9553 (.A1(_00971_),
    .A2(n_9551_o_0),
    .B(n_9552_o_0),
    .Y(n_9553_o_0));
 OAI21xp33_ASAP7_75t_R n_9554 (.A1(n_9417_o_0),
    .A2(n_9546_o_0),
    .B(n_9553_o_0),
    .Y(n_9554_o_0));
 OAI21xp33_ASAP7_75t_R n_9555 (.A1(n_9452_o_0),
    .A2(n_9482_o_0),
    .B(n_9511_o_0),
    .Y(n_9555_o_0));
 NOR2xp33_ASAP7_75t_R n_9556 (.A(n_9435_o_0),
    .B(n_9555_o_0),
    .Y(n_9556_o_0));
 OAI21xp33_ASAP7_75t_R n_9557 (.A1(n_9531_o_0),
    .A2(net53),
    .B(n_9465_o_0),
    .Y(n_9557_o_0));
 AO21x1_ASAP7_75t_R n_9558 (.A1(n_9485_o_0),
    .A2(n_9463_o_0),
    .B(n_9507_o_0),
    .Y(n_9558_o_0));
 AOI21xp33_ASAP7_75t_R n_9559 (.A1(n_9511_o_0),
    .A2(n_9519_o_0),
    .B(n_9531_o_0),
    .Y(n_9559_o_0));
 NAND2xp33_ASAP7_75t_R n_956 (.A(n_859_o_0),
    .B(n_836_o_0),
    .Y(n_956_o_0));
 INVx1_ASAP7_75t_R n_9560 (.A(n_9559_o_0),
    .Y(n_9560_o_0));
 AOI21xp33_ASAP7_75t_R n_9561 (.A1(n_9558_o_0),
    .A2(n_9560_o_0),
    .B(n_9526_o_0),
    .Y(n_9561_o_0));
 OAI21xp33_ASAP7_75t_R n_9562 (.A1(n_9556_o_0),
    .A2(n_9557_o_0),
    .B(n_9561_o_0),
    .Y(n_9562_o_0));
 NAND2xp33_ASAP7_75t_R n_9563 (.A(n_9451_o_0),
    .B(n_9482_o_0),
    .Y(n_9563_o_0));
 NAND3xp33_ASAP7_75t_R n_9564 (.A(n_9531_o_0),
    .B(n_9452_o_0),
    .C(net53),
    .Y(n_9564_o_0));
 OAI211xp5_ASAP7_75t_R n_9565 (.A1(n_9531_o_0),
    .A2(n_9563_o_0),
    .B(n_9564_o_0),
    .C(n_9465_o_0),
    .Y(n_9565_o_0));
 OAI31xp33_ASAP7_75t_R n_9566 (.A1(n_9508_o_0),
    .A2(n_9535_o_0),
    .A3(n_9520_o_0),
    .B(n_9565_o_0),
    .Y(n_9566_o_0));
 INVx1_ASAP7_75t_R n_9567 (.A(n_9422_o_0),
    .Y(n_9567_o_0));
 AOI21xp33_ASAP7_75t_R n_9568 (.A1(n_9526_o_0),
    .A2(n_9566_o_0),
    .B(n_9567_o_0),
    .Y(n_9568_o_0));
 NOR3xp33_ASAP7_75t_R n_9569 (.A(n_9452_o_0),
    .B(net53),
    .C(n_9435_o_0),
    .Y(n_9569_o_0));
 INVx1_ASAP7_75t_R n_957 (.A(n_913_o_0),
    .Y(n_957_o_0));
 INVx1_ASAP7_75t_R n_9570 (.A(n_9569_o_0),
    .Y(n_9570_o_0));
 NAND3xp33_ASAP7_75t_R n_9571 (.A(n_9570_o_0),
    .B(n_9453_o_0),
    .C(n_9558_o_0),
    .Y(n_9571_o_0));
 OAI211xp5_ASAP7_75t_R n_9572 (.A1(n_9435_o_0),
    .A2(n_9452_o_0),
    .B(n_9508_o_0),
    .C(net26),
    .Y(n_9572_o_0));
 AO21x1_ASAP7_75t_R n_9573 (.A1(n_9571_o_0),
    .A2(n_9572_o_0),
    .B(n_9542_o_0),
    .Y(n_9573_o_0));
 INVx1_ASAP7_75t_R n_9574 (.A(n_9453_o_0),
    .Y(n_9574_o_0));
 NOR2xp67_ASAP7_75t_R n_9575 (.A(n_9482_o_0),
    .B(n_9452_o_0),
    .Y(n_9575_o_0));
 NOR2xp33_ASAP7_75t_R n_9576 (.A(n_9435_o_0),
    .B(n_9575_o_0),
    .Y(n_9576_o_0));
 NAND2xp33_ASAP7_75t_R n_9577 (.A(net53),
    .B(n_9531_o_0),
    .Y(n_9577_o_0));
 NAND3xp33_ASAP7_75t_R n_9578 (.A(n_9492_o_0),
    .B(n_9577_o_0),
    .C(n_9465_o_0),
    .Y(n_9578_o_0));
 OAI31xp33_ASAP7_75t_R n_9579 (.A1(n_9508_o_0),
    .A2(n_9574_o_0),
    .A3(n_9576_o_0),
    .B(n_9578_o_0),
    .Y(n_9579_o_0));
 NOR2xp33_ASAP7_75t_R n_958 (.A(n_877_o_0),
    .B(n_945_o_0),
    .Y(n_958_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9580 (.A1(n_9499_o_0),
    .A2(n_1359_o_0),
    .B(n_9500_o_0),
    .C(n_9579_o_0),
    .Y(n_9580_o_0));
 AOI22xp33_ASAP7_75t_R n_9581 (.A1(n_9562_o_0),
    .A2(n_9568_o_0),
    .B1(n_9573_o_0),
    .B2(n_9580_o_0),
    .Y(n_9581_o_0));
 NAND3xp33_ASAP7_75t_R n_9582 (.A(n_9568_o_0),
    .B(n_9562_o_0),
    .C(n_9422_o_0),
    .Y(n_9582_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9583 (.A1(n_9422_o_0),
    .A2(n_9581_o_0),
    .B(n_9582_o_0),
    .C(n_9416_o_1),
    .Y(n_9583_o_0));
 AOI21xp33_ASAP7_75t_R n_9584 (.A1(n_9531_o_0),
    .A2(n_9555_o_0),
    .B(n_9465_o_0),
    .Y(n_9584_o_0));
 AOI21xp33_ASAP7_75t_R n_9585 (.A1(n_9538_o_0),
    .A2(n_9492_o_0),
    .B(n_9558_o_0),
    .Y(n_9585_o_0));
 OAI21xp33_ASAP7_75t_R n_9586 (.A1(n_9584_o_0),
    .A2(n_9585_o_0),
    .B(n_9523_o_0),
    .Y(n_9586_o_0));
 NOR2xp33_ASAP7_75t_R n_9587 (.A(n_9531_o_0),
    .B(n_9558_o_0),
    .Y(n_9587_o_0));
 NAND2xp33_ASAP7_75t_R n_9588 (.A(n_9483_o_0),
    .B(n_9587_o_0),
    .Y(n_9588_o_0));
 AO21x1_ASAP7_75t_R n_9589 (.A1(n_9588_o_0),
    .A2(n_9571_o_0),
    .B(n_9542_o_0),
    .Y(n_9589_o_0));
 OAI21xp33_ASAP7_75t_R n_959 (.A1(n_957_o_0),
    .A2(n_836_o_0),
    .B(n_958_o_0),
    .Y(n_959_o_0));
 AOI21xp33_ASAP7_75t_R n_9590 (.A1(n_9586_o_0),
    .A2(n_9589_o_0),
    .B(n_9544_o_0),
    .Y(n_9590_o_0));
 INVx1_ASAP7_75t_R n_9591 (.A(n_9482_o_0),
    .Y(n_9591_o_0));
 OAI21xp33_ASAP7_75t_R n_9592 (.A1(n_9531_o_0),
    .A2(n_9555_o_0),
    .B(n_9465_o_0),
    .Y(n_9592_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9593 (.A1(n_9531_o_0),
    .A2(n_9591_o_0),
    .B(n_9508_o_0),
    .C(n_9592_o_0),
    .Y(n_9593_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9594 (.A1(n_9435_o_0),
    .A2(net26),
    .B(n_9452_o_0),
    .C(n_9508_o_0),
    .Y(n_9594_o_0));
 INVx1_ASAP7_75t_R n_9595 (.A(n_9483_o_0),
    .Y(n_9595_o_0));
 NAND3xp33_ASAP7_75t_R n_9596 (.A(n_9595_o_0),
    .B(n_9531_o_0),
    .C(n_9508_o_0),
    .Y(n_9596_o_0));
 OAI311xp33_ASAP7_75t_R n_9597 (.A1(n_9558_o_0),
    .A2(n_9531_o_0),
    .A3(n_9451_o_0),
    .B1(n_9526_o_0),
    .C1(n_9596_o_0),
    .Y(n_9597_o_0));
 OAI21xp33_ASAP7_75t_R n_9598 (.A1(n_9594_o_0),
    .A2(n_9597_o_0),
    .B(n_9422_o_0),
    .Y(n_9598_o_0));
 AOI21xp33_ASAP7_75t_R n_9599 (.A1(n_9542_o_0),
    .A2(n_9593_o_0),
    .B(n_9598_o_0),
    .Y(n_9599_o_0));
 AOI31xp33_ASAP7_75t_R n_960 (.A1(n_877_o_0),
    .A2(n_881_o_0),
    .A3(n_860_o_0),
    .B(n_829_o_0),
    .Y(n_960_o_0));
 INVx1_ASAP7_75t_R n_9600 (.A(n_9553_o_0),
    .Y(n_9600_o_0));
 NAND2xp33_ASAP7_75t_R n_9601 (.A(n_9482_o_0),
    .B(n_9452_o_0),
    .Y(n_9601_o_0));
 AOI21xp33_ASAP7_75t_R n_9602 (.A1(n_9452_o_0),
    .A2(net53),
    .B(n_9531_o_0),
    .Y(n_9602_o_0));
 INVx1_ASAP7_75t_R n_9603 (.A(n_9602_o_0),
    .Y(n_9603_o_0));
 OAI31xp33_ASAP7_75t_R n_9604 (.A1(n_9558_o_0),
    .A2(n_9435_o_0),
    .A3(n_9601_o_0),
    .B(n_9603_o_0),
    .Y(n_9604_o_0));
 NAND2xp33_ASAP7_75t_R n_9605 (.A(n_9508_o_0),
    .B(n_9604_o_0),
    .Y(n_9605_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9606 (.A1(n_9435_o_0),
    .A2(net22),
    .B(n_9490_o_0),
    .C(n_9501_o_0),
    .Y(n_9606_o_0));
 NOR2xp33_ASAP7_75t_R n_9607 (.A(n_9531_o_0),
    .B(n_9563_o_0),
    .Y(n_9607_o_0));
 NOR3xp33_ASAP7_75t_R n_9608 (.A(n_9607_o_0),
    .B(n_9505_o_0),
    .C(n_9508_o_0),
    .Y(n_9608_o_0));
 NOR2xp33_ASAP7_75t_R n_9609 (.A(n_9482_o_0),
    .B(n_9435_o_0),
    .Y(n_9609_o_0));
 OA211x2_ASAP7_75t_R n_961 (.A1(n_956_o_0),
    .A2(n_878_o_0),
    .B(n_959_o_0),
    .C(n_960_o_0),
    .Y(n_961_o_0));
 OAI21xp33_ASAP7_75t_R n_9610 (.A1(n_9609_o_0),
    .A2(n_9592_o_0),
    .B(n_9501_o_0),
    .Y(n_9610_o_0));
 OAI21xp33_ASAP7_75t_R n_9611 (.A1(n_9608_o_0),
    .A2(n_9610_o_0),
    .B(n_9567_o_0),
    .Y(n_9611_o_0));
 NOR3xp33_ASAP7_75t_R n_9612 (.A(n_9601_o_0),
    .B(n_9465_o_0),
    .C(n_9435_o_0),
    .Y(n_9612_o_0));
 OAI31xp33_ASAP7_75t_R n_9613 (.A1(n_9452_o_0),
    .A2(n_9591_o_0),
    .A3(n_9531_o_0),
    .B(n_9465_o_0),
    .Y(n_9613_o_0));
 AOI21xp33_ASAP7_75t_R n_9614 (.A1(n_9531_o_0),
    .A2(net22),
    .B(n_9613_o_0),
    .Y(n_9614_o_0));
 OAI31xp33_ASAP7_75t_R n_9615 (.A1(n_9451_o_0),
    .A2(n_9435_o_0),
    .A3(net53),
    .B(n_9558_o_0),
    .Y(n_9615_o_0));
 AOI21xp33_ASAP7_75t_R n_9616 (.A1(n_9451_o_0),
    .A2(n_9482_o_0),
    .B(n_9531_o_0),
    .Y(n_9616_o_0));
 OAI321xp33_ASAP7_75t_R n_9617 (.A1(n_9558_o_0),
    .A2(n_9435_o_0),
    .A3(n_9601_o_0),
    .B1(n_9615_o_0),
    .B2(n_9616_o_0),
    .C(n_9501_o_0),
    .Y(n_9617_o_0));
 OAI31xp33_ASAP7_75t_R n_9618 (.A1(n_9501_o_0),
    .A2(n_9612_o_0),
    .A3(n_9614_o_0),
    .B(n_9617_o_0),
    .Y(n_9618_o_0));
 OAI21xp33_ASAP7_75t_R n_9619 (.A1(n_9415_o_0),
    .A2(n_1422_o_0),
    .B(n_9416_o_0),
    .Y(n_9619_o_0));
 AOI211xp5_ASAP7_75t_R n_962 (.A1(n_951_o_0),
    .A2(n_955_o_0),
    .B(n_961_o_0),
    .C(n_904_o_0),
    .Y(n_962_o_0));
 OA21x2_ASAP7_75t_R n_9620 (.A1(n_9618_o_0),
    .A2(n_9567_o_0),
    .B(n_9619_o_0),
    .Y(n_9620_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9621 (.A1(n_9605_o_0),
    .A2(n_9606_o_0),
    .B(n_9611_o_0),
    .C(n_9620_o_0),
    .Y(n_9621_o_0));
 OAI311xp33_ASAP7_75t_R n_9622 (.A1(n_9416_o_1),
    .A2(n_9590_o_0),
    .A3(n_9599_o_0),
    .B1(n_9600_o_0),
    .C1(n_9621_o_0),
    .Y(n_9622_o_0));
 OAI21xp33_ASAP7_75t_R n_9623 (.A1(n_9554_o_0),
    .A2(n_9583_o_0),
    .B(n_9622_o_0),
    .Y(n_9623_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9624 (.A1(n_9519_o_0),
    .A2(n_9511_o_0),
    .B(n_9531_o_0),
    .C(n_9490_o_0),
    .Y(n_9624_o_0));
 NOR2xp33_ASAP7_75t_R n_9625 (.A(n_9435_o_0),
    .B(n_9575_o_0),
    .Y(n_9625_o_0));
 OAI211xp5_ASAP7_75t_R n_9626 (.A1(n_9624_o_0),
    .A2(n_9625_o_0),
    .B(n_9596_o_0),
    .C(n_9526_o_0),
    .Y(n_9626_o_0));
 NAND2xp33_ASAP7_75t_R n_9627 (.A(n_9435_o_0),
    .B(n_9591_o_0),
    .Y(n_9627_o_0));
 AOI21xp33_ASAP7_75t_R n_9628 (.A1(n_9558_o_0),
    .A2(n_9627_o_0),
    .B(n_9501_o_0),
    .Y(n_9628_o_0));
 OAI21xp33_ASAP7_75t_R n_9629 (.A1(n_9558_o_0),
    .A2(n_9577_o_0),
    .B(n_9628_o_0),
    .Y(n_9629_o_0));
 AOI211xp5_ASAP7_75t_R n_963 (.A1(n_904_o_0),
    .A2(n_948_o_0),
    .B(n_962_o_0),
    .C(n_930_o_0),
    .Y(n_963_o_0));
 AO21x1_ASAP7_75t_R n_9630 (.A1(n_9626_o_0),
    .A2(n_9629_o_0),
    .B(n_9416_o_1),
    .Y(n_9630_o_0));
 NOR2xp33_ASAP7_75t_R n_9631 (.A(n_1422_o_0),
    .B(n_9415_o_0),
    .Y(n_9631_o_0));
 AOI21xp33_ASAP7_75t_R n_9632 (.A1(n_1422_o_0),
    .A2(n_9415_o_0),
    .B(n_9631_o_0),
    .Y(n_9632_o_0));
 NOR2xp33_ASAP7_75t_R n_9633 (.A(n_9632_o_0),
    .B(n_9523_o_0),
    .Y(n_9633_o_0));
 AOI211xp5_ASAP7_75t_R n_9634 (.A1(n_9452_o_0),
    .A2(net26),
    .B(n_9609_o_0),
    .C(n_9490_o_0),
    .Y(n_9634_o_0));
 AOI31xp33_ASAP7_75t_R n_9635 (.A1(n_9558_o_0),
    .A2(n_9595_o_0),
    .A3(n_9435_o_0),
    .B(n_9634_o_0),
    .Y(n_9635_o_0));
 AOI21xp33_ASAP7_75t_R n_9636 (.A1(n_9451_o_0),
    .A2(n_9435_o_0),
    .B(n_9490_o_0),
    .Y(n_9636_o_0));
 OAI21xp33_ASAP7_75t_R n_9637 (.A1(n_9451_o_0),
    .A2(net53),
    .B(n_9531_o_0),
    .Y(n_9637_o_0));
 AOI211xp5_ASAP7_75t_R n_9638 (.A1(n_9636_o_0),
    .A2(n_9637_o_0),
    .B(n_9632_o_0),
    .C(n_9501_o_0),
    .Y(n_9638_o_0));
 OAI31xp33_ASAP7_75t_R n_9639 (.A1(n_9508_o_0),
    .A2(n_9574_o_0),
    .A3(net85),
    .B(n_9638_o_0),
    .Y(n_9639_o_0));
 INVx1_ASAP7_75t_R n_964 (.A(_00979_),
    .Y(n_964_o_0));
 INVx1_ASAP7_75t_R n_9640 (.A(n_9639_o_0),
    .Y(n_9640_o_0));
 AOI21xp33_ASAP7_75t_R n_9641 (.A1(n_9633_o_0),
    .A2(n_9635_o_0),
    .B(n_9640_o_0),
    .Y(n_9641_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9642 (.A1(net22),
    .A2(n_9587_o_0),
    .B(n_9630_o_0),
    .C(n_9641_o_0),
    .Y(n_9642_o_0));
 AOI21xp33_ASAP7_75t_R n_9643 (.A1(n_9482_o_0),
    .A2(n_9452_o_0),
    .B(n_9435_o_0),
    .Y(n_9643_o_0));
 INVx1_ASAP7_75t_R n_9644 (.A(n_9643_o_0),
    .Y(n_9644_o_0));
 AOI21xp33_ASAP7_75t_R n_9645 (.A1(n_9636_o_0),
    .A2(n_9644_o_0),
    .B(n_9526_o_0),
    .Y(n_9645_o_0));
 OAI31xp33_ASAP7_75t_R n_9646 (.A1(n_9508_o_0),
    .A2(n_9493_o_0),
    .A3(net85),
    .B(n_9645_o_0),
    .Y(n_9646_o_0));
 NOR2xp33_ASAP7_75t_R n_9647 (.A(n_9508_o_0),
    .B(n_9505_o_0),
    .Y(n_9647_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9648 (.A1(n_9452_o_0),
    .A2(net26),
    .B(n_9647_o_0),
    .C(n_9542_o_0),
    .Y(n_9648_o_0));
 OAI31xp33_ASAP7_75t_R n_9649 (.A1(n_9490_o_0),
    .A2(n_9559_o_0),
    .A3(n_9529_o_0),
    .B(n_9648_o_0),
    .Y(n_9649_o_0));
 XNOR2xp5_ASAP7_75t_R n_965 (.A(_00445_),
    .B(_00883_),
    .Y(n_965_o_0));
 NAND3xp33_ASAP7_75t_R n_9650 (.A(n_9646_o_0),
    .B(n_9649_o_0),
    .C(n_9417_o_0),
    .Y(n_9650_o_0));
 NAND2xp33_ASAP7_75t_R n_9651 (.A(n_9451_o_0),
    .B(n_9591_o_0),
    .Y(n_9651_o_0));
 NOR2xp33_ASAP7_75t_R n_9652 (.A(n_9435_o_0),
    .B(n_9591_o_0),
    .Y(n_9652_o_0));
 NOR3xp33_ASAP7_75t_R n_9653 (.A(n_9510_o_0),
    .B(n_9652_o_0),
    .C(n_9508_o_0),
    .Y(n_9653_o_0));
 AOI31xp33_ASAP7_75t_R n_9654 (.A1(n_9531_o_0),
    .A2(n_9651_o_0),
    .A3(n_9465_o_0),
    .B(n_9653_o_0),
    .Y(n_9654_o_0));
 AOI21xp33_ASAP7_75t_R n_9655 (.A1(n_9435_o_0),
    .A2(n_9575_o_0),
    .B(n_9508_o_0),
    .Y(n_9655_o_0));
 OAI21xp33_ASAP7_75t_R n_9656 (.A1(n_9435_o_0),
    .A2(n_9555_o_0),
    .B(n_9655_o_0),
    .Y(n_9656_o_0));
 OAI31xp33_ASAP7_75t_R n_9657 (.A1(n_9435_o_0),
    .A2(n_9490_o_0),
    .A3(n_9595_o_0),
    .B(n_9656_o_0),
    .Y(n_9657_o_0));
 AOI21xp33_ASAP7_75t_R n_9658 (.A1(n_9526_o_0),
    .A2(n_9657_o_0),
    .B(n_9417_o_0),
    .Y(n_9658_o_0));
 OAI21xp33_ASAP7_75t_R n_9659 (.A1(n_9501_o_0),
    .A2(n_9654_o_0),
    .B(n_9658_o_0),
    .Y(n_9659_o_0));
 XNOR2xp5_ASAP7_75t_R n_966 (.A(_00915_),
    .B(n_965_o_0),
    .Y(n_966_o_0));
 INVx1_ASAP7_75t_R n_9660 (.A(n_9544_o_0),
    .Y(n_9660_o_0));
 XNOR2xp5_ASAP7_75t_R n_9661 (.A(_00971_),
    .B(n_9551_o_0),
    .Y(n_9661_o_0));
 AOI31xp33_ASAP7_75t_R n_9662 (.A1(n_9650_o_0),
    .A2(n_9659_o_0),
    .A3(n_9660_o_0),
    .B(n_9661_o_0),
    .Y(n_9662_o_0));
 OAI21xp33_ASAP7_75t_R n_9663 (.A1(n_9435_o_0),
    .A2(n_9575_o_0),
    .B(n_9465_o_0),
    .Y(n_9663_o_0));
 OAI21xp33_ASAP7_75t_R n_9664 (.A1(n_9602_o_0),
    .A2(n_9663_o_0),
    .B(n_9632_o_0),
    .Y(n_9664_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9665 (.A1(n_9555_o_0),
    .A2(n_9435_o_0),
    .B(n_9655_o_0),
    .C(n_9664_o_0),
    .Y(n_9665_o_0));
 AOI31xp33_ASAP7_75t_R n_9666 (.A1(n_9511_o_0),
    .A2(n_9519_o_0),
    .A3(n_9435_o_0),
    .B(n_9508_o_0),
    .Y(n_9666_o_0));
 AOI21xp33_ASAP7_75t_R n_9667 (.A1(n_9644_o_0),
    .A2(n_9666_o_0),
    .B(n_9636_o_0),
    .Y(n_9667_o_0));
 NOR3xp33_ASAP7_75t_R n_9668 (.A(n_9558_o_0),
    .B(n_9601_o_0),
    .C(n_9435_o_0),
    .Y(n_9668_o_0));
 NOR3xp33_ASAP7_75t_R n_9669 (.A(n_9667_o_0),
    .B(n_9632_o_0),
    .C(n_9668_o_0),
    .Y(n_9669_o_0));
 XNOR2xp5_ASAP7_75t_R n_967 (.A(_00947_),
    .B(n_966_o_0),
    .Y(n_967_o_0));
 OAI32xp33_ASAP7_75t_R n_9670 (.A1(n_9569_o_0),
    .A2(n_9574_o_0),
    .A3(n_9490_o_0),
    .B1(n_9520_o_0),
    .B2(n_9508_o_0),
    .Y(n_9670_o_0));
 NAND2xp33_ASAP7_75t_R n_9671 (.A(n_9482_o_0),
    .B(n_9435_o_0),
    .Y(n_9671_o_0));
 NAND3xp33_ASAP7_75t_R n_9672 (.A(n_9558_o_0),
    .B(n_9671_o_0),
    .C(n_9637_o_0),
    .Y(n_9672_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9673 (.A1(n_9490_o_0),
    .A2(n_9535_o_0),
    .B(n_9672_o_0),
    .C(n_9529_o_0),
    .Y(n_9673_o_0));
 OAI221xp5_ASAP7_75t_R n_9674 (.A1(n_9619_o_0),
    .A2(n_9670_o_0),
    .B1(n_9417_o_0),
    .B2(n_9673_o_0),
    .C(n_9526_o_0),
    .Y(n_9674_o_0));
 OAI31xp33_ASAP7_75t_R n_9675 (.A1(n_9501_o_0),
    .A2(n_9665_o_0),
    .A3(n_9669_o_0),
    .B(n_9674_o_0),
    .Y(n_9675_o_0));
 OAI21xp33_ASAP7_75t_R n_9676 (.A1(n_9569_o_0),
    .A2(n_9613_o_0),
    .B(n_9501_o_0),
    .Y(n_9676_o_0));
 INVx1_ASAP7_75t_R n_9677 (.A(n_9676_o_0),
    .Y(n_9677_o_0));
 NAND2xp33_ASAP7_75t_R n_9678 (.A(net26),
    .B(n_9435_o_0),
    .Y(n_9678_o_0));
 NAND3xp33_ASAP7_75t_R n_9679 (.A(n_9417_o_0),
    .B(n_9558_o_0),
    .C(n_9678_o_0),
    .Y(n_9679_o_0));
 INVx1_ASAP7_75t_R n_968 (.A(n_967_o_0),
    .Y(n_968_o_0));
 NOR2xp33_ASAP7_75t_R n_9680 (.A(n_9490_o_0),
    .B(n_9505_o_0),
    .Y(n_9680_o_0));
 INVx1_ASAP7_75t_R n_9681 (.A(n_9680_o_0),
    .Y(n_9681_o_0));
 AOI21xp33_ASAP7_75t_R n_9682 (.A1(n_9435_o_0),
    .A2(n_9483_o_0),
    .B(n_9508_o_0),
    .Y(n_9682_o_0));
 AOI21xp33_ASAP7_75t_R n_9683 (.A1(n_9682_o_0),
    .A2(n_9570_o_0),
    .B(n_9417_o_0),
    .Y(n_9683_o_0));
 OAI21xp33_ASAP7_75t_R n_9684 (.A1(n_9681_o_0),
    .A2(n_9535_o_0),
    .B(n_9683_o_0),
    .Y(n_9684_o_0));
 AOI31xp33_ASAP7_75t_R n_9685 (.A1(n_9558_o_0),
    .A2(n_9671_o_0),
    .A3(n_9637_o_0),
    .B(n_9619_o_0),
    .Y(n_9685_o_0));
 OAI21xp33_ASAP7_75t_R n_9686 (.A1(n_9557_o_0),
    .A2(n_9529_o_0),
    .B(n_9685_o_0),
    .Y(n_9686_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9687 (.A1(n_9684_o_0),
    .A2(n_9686_o_0),
    .B(n_9526_o_0),
    .C(n_9544_o_0),
    .Y(n_9687_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9688 (.A1(n_9677_o_0),
    .A2(n_9679_o_0),
    .B(n_9687_o_0),
    .C(n_9661_o_0),
    .Y(n_9688_o_0));
 AOI21xp33_ASAP7_75t_R n_9689 (.A1(n_9567_o_0),
    .A2(n_9675_o_0),
    .B(n_9688_o_0),
    .Y(n_9689_o_0));
 NOR2xp33_ASAP7_75t_R n_969 (.A(n_964_o_0),
    .B(n_968_o_0),
    .Y(n_969_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9690 (.A1(n_9567_o_0),
    .A2(n_9642_o_0),
    .B(n_9662_o_0),
    .C(n_9689_o_0),
    .Y(n_9690_o_0));
 AOI21xp33_ASAP7_75t_R n_9691 (.A1(n_9435_o_0),
    .A2(n_9483_o_0),
    .B(n_9508_o_0),
    .Y(n_9691_o_0));
 OAI21xp33_ASAP7_75t_R n_9692 (.A1(n_9531_o_0),
    .A2(n_9651_o_0),
    .B(n_9508_o_0),
    .Y(n_9692_o_0));
 OAI21xp33_ASAP7_75t_R n_9693 (.A1(n_9539_o_0),
    .A2(n_9692_o_0),
    .B(n_9523_o_0),
    .Y(n_9693_o_0));
 AOI21xp33_ASAP7_75t_R n_9694 (.A1(n_9691_o_0),
    .A2(n_9532_o_0),
    .B(n_9693_o_0),
    .Y(n_9694_o_0));
 NAND2xp33_ASAP7_75t_R n_9695 (.A(net26),
    .B(n_9531_o_0),
    .Y(n_9695_o_0));
 AOI21xp33_ASAP7_75t_R n_9696 (.A1(n_9435_o_0),
    .A2(n_9595_o_0),
    .B(n_9465_o_0),
    .Y(n_9696_o_0));
 AOI21xp33_ASAP7_75t_R n_9697 (.A1(n_9695_o_0),
    .A2(n_9696_o_0),
    .B(n_9585_o_0),
    .Y(n_9697_o_0));
 OAI21xp33_ASAP7_75t_R n_9698 (.A1(n_9542_o_0),
    .A2(n_9697_o_0),
    .B(n_9417_o_0),
    .Y(n_9698_o_0));
 NAND2xp33_ASAP7_75t_R n_9699 (.A(n_9671_o_0),
    .B(n_9558_o_0),
    .Y(n_9699_o_0));
 AOI211xp5_ASAP7_75t_R n_970 (.A1(n_964_o_0),
    .A2(n_968_o_0),
    .B(n_969_o_0),
    .C(ld),
    .Y(n_970_o_0));
 INVx1_ASAP7_75t_R n_9700 (.A(n_9692_o_0),
    .Y(n_9700_o_0));
 AOI21xp33_ASAP7_75t_R n_9701 (.A1(n_9532_o_0),
    .A2(n_9700_o_0),
    .B(n_9526_o_0),
    .Y(n_9701_o_0));
 OAI21xp33_ASAP7_75t_R n_9702 (.A1(n_9699_o_0),
    .A2(n_9539_o_0),
    .B(n_9701_o_0),
    .Y(n_9702_o_0));
 INVx1_ASAP7_75t_R n_9703 (.A(n_9520_o_0),
    .Y(n_9703_o_0));
 NAND2xp33_ASAP7_75t_R n_9704 (.A(n_9666_o_0),
    .B(n_9703_o_0),
    .Y(n_9704_o_0));
 OAI31xp33_ASAP7_75t_R n_9705 (.A1(n_9490_o_0),
    .A2(n_9505_o_0),
    .A3(n_9616_o_0),
    .B(n_9704_o_0),
    .Y(n_9705_o_0));
 AOI21xp33_ASAP7_75t_R n_9706 (.A1(n_9526_o_0),
    .A2(n_9705_o_0),
    .B(n_9417_o_0),
    .Y(n_9706_o_0));
 AOI21xp33_ASAP7_75t_R n_9707 (.A1(n_9702_o_0),
    .A2(n_9706_o_0),
    .B(n_9544_o_0),
    .Y(n_9707_o_0));
 OAI21xp33_ASAP7_75t_R n_9708 (.A1(n_9694_o_0),
    .A2(n_9698_o_0),
    .B(n_9707_o_0),
    .Y(n_9708_o_0));
 OA21x2_ASAP7_75t_R n_9709 (.A1(n_9435_o_0),
    .A2(n_9483_o_0),
    .B(n_9691_o_0),
    .Y(n_9709_o_0));
 AOI21xp33_ASAP7_75t_R n_971 (.A1(key[23]),
    .A2(ld),
    .B(n_970_o_0),
    .Y(n_971_o_0));
 INVx1_ASAP7_75t_R n_9710 (.A(n_9637_o_0),
    .Y(n_9710_o_0));
 OAI21xp33_ASAP7_75t_R n_9711 (.A1(n_9435_o_0),
    .A2(net26),
    .B(n_9682_o_0),
    .Y(n_9711_o_0));
 OAI31xp33_ASAP7_75t_R n_9712 (.A1(n_9490_o_0),
    .A2(n_9510_o_0),
    .A3(n_9710_o_0),
    .B(n_9711_o_0),
    .Y(n_9712_o_0));
 AOI21xp33_ASAP7_75t_R n_9713 (.A1(n_9542_o_0),
    .A2(n_9712_o_0),
    .B(n_9416_o_1),
    .Y(n_9713_o_0));
 OAI21xp33_ASAP7_75t_R n_9714 (.A1(n_9610_o_0),
    .A2(n_9709_o_0),
    .B(n_9713_o_0),
    .Y(n_9714_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9715 (.A1(n_9435_o_0),
    .A2(n_9575_o_0),
    .B(n_9655_o_0),
    .C(n_9504_o_0),
    .Y(n_9715_o_0));
 OAI211xp5_ASAP7_75t_R n_9716 (.A1(n_9555_o_0),
    .A2(n_9435_o_0),
    .B(n_9465_o_0),
    .C(n_9671_o_0),
    .Y(n_9716_o_0));
 OAI211xp5_ASAP7_75t_R n_9717 (.A1(n_9601_o_0),
    .A2(n_9531_o_0),
    .B(n_9558_o_0),
    .C(n_9532_o_0),
    .Y(n_9717_o_0));
 AOI31xp33_ASAP7_75t_R n_9718 (.A1(n_9523_o_0),
    .A2(n_9716_o_0),
    .A3(n_9717_o_0),
    .B(n_9632_o_0),
    .Y(n_9718_o_0));
 OAI21xp33_ASAP7_75t_R n_9719 (.A1(n_9542_o_0),
    .A2(n_9715_o_0),
    .B(n_9718_o_0),
    .Y(n_9719_o_0));
 INVx1_ASAP7_75t_R n_972 (.A(n_971_o_0),
    .Y(n_972_o_0));
 NAND3xp33_ASAP7_75t_R n_9720 (.A(n_9714_o_0),
    .B(n_9719_o_0),
    .C(n_9422_o_0),
    .Y(n_9720_o_0));
 INVx1_ASAP7_75t_R n_9721 (.A(n_9661_o_0),
    .Y(n_9721_o_0));
 AOI21xp33_ASAP7_75t_R n_9722 (.A1(n_9481_o_0),
    .A2(n_9518_o_0),
    .B(n_9451_o_0),
    .Y(n_9722_o_0));
 AOI211xp5_ASAP7_75t_R n_9723 (.A1(_00964_),
    .A2(n_9444_o_0),
    .B(net53),
    .C(n_9450_o_0),
    .Y(n_9723_o_0));
 OAI21xp33_ASAP7_75t_R n_9724 (.A1(n_9452_o_0),
    .A2(n_9591_o_0),
    .B(n_9531_o_0),
    .Y(n_9724_o_0));
 OAI311xp33_ASAP7_75t_R n_9725 (.A1(n_9531_o_0),
    .A2(n_9722_o_0),
    .A3(n_9723_o_0),
    .B1(n_9558_o_0),
    .C1(n_9724_o_0),
    .Y(n_9725_o_0));
 OAI31xp33_ASAP7_75t_R n_9726 (.A1(n_9490_o_0),
    .A2(n_9602_o_0),
    .A3(n_9609_o_0),
    .B(n_9725_o_0),
    .Y(n_9726_o_0));
 AOI21xp33_ASAP7_75t_R n_9727 (.A1(n_9542_o_0),
    .A2(n_9726_o_0),
    .B(n_9619_o_0),
    .Y(n_9727_o_0));
 AOI311xp33_ASAP7_75t_R n_9728 (.A1(net89),
    .A2(n_9519_o_0),
    .A3(n_9435_o_0),
    .B(n_9490_o_0),
    .C(n_9609_o_0),
    .Y(n_9728_o_0));
 AOI31xp33_ASAP7_75t_R n_9729 (.A1(n_9558_o_0),
    .A2(n_9671_o_0),
    .A3(n_9506_o_0),
    .B(n_9728_o_0),
    .Y(n_9729_o_0));
 NAND3xp33_ASAP7_75t_R n_973 (.A(n_910_o_0),
    .B(n_865_o_0),
    .C(n_878_o_0),
    .Y(n_973_o_0));
 AOI21xp33_ASAP7_75t_R n_9730 (.A1(n_9542_o_0),
    .A2(n_9729_o_0),
    .B(n_9632_o_0),
    .Y(n_9730_o_0));
 INVx1_ASAP7_75t_R n_9731 (.A(n_9678_o_0),
    .Y(n_9731_o_0));
 OAI211xp5_ASAP7_75t_R n_9732 (.A1(net26),
    .A2(n_9435_o_0),
    .B(n_9558_o_0),
    .C(n_9527_o_0),
    .Y(n_9732_o_0));
 OA21x2_ASAP7_75t_R n_9733 (.A1(n_9490_o_0),
    .A2(n_9731_o_0),
    .B(n_9732_o_0),
    .Y(n_9733_o_0));
 NOR3xp33_ASAP7_75t_R n_9734 (.A(n_9435_o_0),
    .B(net26),
    .C(n_9451_o_0),
    .Y(n_9734_o_0));
 NAND2xp33_ASAP7_75t_R n_9735 (.A(n_9531_o_0),
    .B(n_9591_o_0),
    .Y(n_9735_o_0));
 OAI22xp33_ASAP7_75t_R n_9736 (.A1(n_9624_o_0),
    .A2(n_9734_o_0),
    .B1(n_9558_o_0),
    .B2(n_9735_o_0),
    .Y(n_9736_o_0));
 AOI21xp33_ASAP7_75t_R n_9737 (.A1(n_9619_o_0),
    .A2(n_9736_o_0),
    .B(n_9542_o_0),
    .Y(n_9737_o_0));
 OAI21xp33_ASAP7_75t_R n_9738 (.A1(n_9416_o_1),
    .A2(n_9733_o_0),
    .B(n_9737_o_0),
    .Y(n_9738_o_0));
 OAI21xp33_ASAP7_75t_R n_9739 (.A1(n_9727_o_0),
    .A2(n_9730_o_0),
    .B(n_9738_o_0),
    .Y(n_9739_o_0));
 OAI31xp33_ASAP7_75t_R n_974 (.A1(n_878_o_0),
    .A2(n_892_o_0),
    .A3(n_952_o_0),
    .B(n_973_o_0),
    .Y(n_974_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9740 (.A1(n_9644_o_0),
    .A2(net22),
    .B(n_9655_o_0),
    .C(n_9417_o_0),
    .Y(n_9740_o_0));
 OAI21xp33_ASAP7_75t_R n_9741 (.A1(n_9569_o_0),
    .A2(n_9613_o_0),
    .B(n_9740_o_0),
    .Y(n_9741_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9742 (.A1(net26),
    .A2(n_9435_o_0),
    .B(n_9682_o_0),
    .C(n_9619_o_0),
    .Y(n_9742_o_0));
 OAI21xp33_ASAP7_75t_R n_9743 (.A1(n_9627_o_0),
    .A2(n_9490_o_0),
    .B(n_9742_o_0),
    .Y(n_9743_o_0));
 OAI31xp33_ASAP7_75t_R n_9744 (.A1(n_9722_o_0),
    .A2(n_9723_o_0),
    .A3(n_9465_o_0),
    .B(n_9531_o_0),
    .Y(n_9744_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9745 (.A1(n_9490_o_0),
    .A2(net22),
    .B(n_9531_o_0),
    .C(n_9744_o_0),
    .Y(n_9745_o_0));
 AOI21xp33_ASAP7_75t_R n_9746 (.A1(n_9508_o_0),
    .A2(n_9643_o_0),
    .B(n_9632_o_0),
    .Y(n_9746_o_0));
 AOI211xp5_ASAP7_75t_R n_9747 (.A1(n_9558_o_0),
    .A2(n_9735_o_0),
    .B(n_9504_o_0),
    .C(n_9619_o_0),
    .Y(n_9747_o_0));
 AOI211xp5_ASAP7_75t_R n_9748 (.A1(n_9745_o_0),
    .A2(n_9746_o_0),
    .B(n_9542_o_0),
    .C(n_9747_o_0),
    .Y(n_9748_o_0));
 AOI31xp33_ASAP7_75t_R n_9749 (.A1(n_9542_o_0),
    .A2(n_9741_o_0),
    .A3(n_9743_o_0),
    .B(n_9748_o_0),
    .Y(n_9749_o_0));
 NAND3xp33_ASAP7_75t_R n_975 (.A(n_860_o_0),
    .B(n_881_o_0),
    .C(n_877_o_0),
    .Y(n_975_o_0));
 OAI22xp33_ASAP7_75t_R n_9750 (.A1(n_9739_o_0),
    .A2(n_9422_o_0),
    .B1(n_9660_o_0),
    .B2(n_9749_o_0),
    .Y(n_9750_o_0));
 NAND2xp33_ASAP7_75t_R n_9751 (.A(n_9721_o_0),
    .B(n_9750_o_0),
    .Y(n_9751_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9752 (.A1(n_9708_o_0),
    .A2(n_9720_o_0),
    .B(n_9721_o_0),
    .C(n_9751_o_0),
    .Y(n_9752_o_0));
 NOR2xp33_ASAP7_75t_R n_9753 (.A(n_9490_o_0),
    .B(n_9520_o_0),
    .Y(n_9753_o_0));
 NAND3xp33_ASAP7_75t_R n_9754 (.A(n_9531_o_0),
    .B(net53),
    .C(n_9451_o_0),
    .Y(n_9754_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9755 (.A1(n_9451_o_0),
    .A2(n_9531_o_0),
    .B(n_9754_o_0),
    .C(n_9508_o_0),
    .Y(n_9755_o_0));
 AOI21xp33_ASAP7_75t_R n_9756 (.A1(n_9509_o_0),
    .A2(n_9753_o_0),
    .B(n_9755_o_0),
    .Y(n_9756_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9757 (.A1(n_9435_o_0),
    .A2(net26),
    .B(n_9452_o_0),
    .C(n_9508_o_0),
    .Y(n_9757_o_0));
 OAI21xp33_ASAP7_75t_R n_9758 (.A1(n_9634_o_0),
    .A2(n_9757_o_0),
    .B(n_9526_o_0),
    .Y(n_9758_o_0));
 OAI21xp33_ASAP7_75t_R n_9759 (.A1(n_9501_o_0),
    .A2(n_9756_o_0),
    .B(n_9758_o_0),
    .Y(n_9759_o_0));
 AOI21xp33_ASAP7_75t_R n_976 (.A1(n_975_o_0),
    .A2(n_916_o_0),
    .B(n_878_o_0),
    .Y(n_976_o_0));
 NOR2xp33_ASAP7_75t_R n_9760 (.A(n_9529_o_0),
    .B(n_9692_o_0),
    .Y(n_9760_o_0));
 INVx1_ASAP7_75t_R n_9761 (.A(n_9616_o_0),
    .Y(n_9761_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9762 (.A1(net53),
    .A2(n_9451_o_0),
    .B(n_9643_o_0),
    .C(n_9508_o_0),
    .Y(n_9762_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9763 (.A1(n_9761_o_0),
    .A2(n_9762_o_0),
    .B(n_9676_o_0),
    .C(n_9417_o_0),
    .Y(n_9763_o_0));
 AOI21xp33_ASAP7_75t_R n_9764 (.A1(n_9523_o_0),
    .A2(n_9760_o_0),
    .B(n_9763_o_0),
    .Y(n_9764_o_0));
 AOI21xp33_ASAP7_75t_R n_9765 (.A1(n_9619_o_0),
    .A2(n_9759_o_0),
    .B(n_9764_o_0),
    .Y(n_9765_o_0));
 NAND2xp33_ASAP7_75t_R n_9766 (.A(n_9451_o_0),
    .B(n_9435_o_0),
    .Y(n_9766_o_0));
 AO21x1_ASAP7_75t_R n_9767 (.A1(n_9527_o_0),
    .A2(n_9766_o_0),
    .B(n_9558_o_0),
    .Y(n_9767_o_0));
 INVx1_ASAP7_75t_R n_9768 (.A(n_9682_o_0),
    .Y(n_9768_o_0));
 AOI21xp33_ASAP7_75t_R n_9769 (.A1(n_9767_o_0),
    .A2(n_9768_o_0),
    .B(n_9523_o_0),
    .Y(n_9769_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_977 (.A1(n_941_o_0),
    .A2(n_878_o_0),
    .B(n_976_o_0),
    .C(net42),
    .Y(n_977_o_0));
 AOI311xp33_ASAP7_75t_R n_9770 (.A1(n_9531_o_0),
    .A2(net89),
    .A3(n_9519_o_0),
    .B(n_9490_o_0),
    .C(n_9616_o_0),
    .Y(n_9770_o_0));
 AOI31xp33_ASAP7_75t_R n_9771 (.A1(n_9558_o_0),
    .A2(n_9577_o_0),
    .A3(n_9509_o_0),
    .B(n_9770_o_0),
    .Y(n_9771_o_0));
 OAI21xp33_ASAP7_75t_R n_9772 (.A1(n_9501_o_0),
    .A2(n_9771_o_0),
    .B(n_9632_o_0),
    .Y(n_9772_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9773 (.A1(n_9527_o_0),
    .A2(n_9532_o_0),
    .B(n_9465_o_0),
    .C(n_9523_o_0),
    .Y(n_9773_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9774 (.A1(n_9519_o_0),
    .A2(net89),
    .B(n_9435_o_0),
    .C(n_9508_o_0),
    .Y(n_9774_o_0));
 AOI21xp33_ASAP7_75t_R n_9775 (.A1(n_9435_o_0),
    .A2(n_9563_o_0),
    .B(n_9774_o_0),
    .Y(n_9775_o_0));
 OAI311xp33_ASAP7_75t_R n_9776 (.A1(n_9531_o_0),
    .A2(net26),
    .A3(n_9451_o_0),
    .B1(n_9538_o_0),
    .C1(n_9558_o_0),
    .Y(n_9776_o_0));
 OAI31xp33_ASAP7_75t_R n_9777 (.A1(n_9490_o_0),
    .A2(n_9569_o_0),
    .A3(n_9559_o_0),
    .B(n_9776_o_0),
    .Y(n_9777_o_0));
 AOI21xp33_ASAP7_75t_R n_9778 (.A1(n_9526_o_0),
    .A2(n_9777_o_0),
    .B(n_9417_o_0),
    .Y(n_9778_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9779 (.A1(n_9773_o_0),
    .A2(n_9775_o_0),
    .B(n_9778_o_0),
    .C(n_9661_o_0),
    .Y(n_9779_o_0));
 OAI211xp5_ASAP7_75t_R n_978 (.A1(net16),
    .A2(n_974_o_0),
    .B(n_977_o_0),
    .C(n_904_o_0),
    .Y(n_978_o_0));
 OAI21xp33_ASAP7_75t_R n_9780 (.A1(n_9769_o_0),
    .A2(n_9772_o_0),
    .B(n_9779_o_0),
    .Y(n_9780_o_0));
 OA21x2_ASAP7_75t_R n_9781 (.A1(n_9765_o_0),
    .A2(n_9600_o_0),
    .B(n_9780_o_0),
    .Y(n_9781_o_0));
 OAI21xp33_ASAP7_75t_R n_9782 (.A1(n_9435_o_0),
    .A2(n_9575_o_0),
    .B(n_9696_o_0),
    .Y(n_9782_o_0));
 AOI21xp33_ASAP7_75t_R n_9783 (.A1(n_9490_o_0),
    .A2(n_9559_o_0),
    .B(n_9416_o_1),
    .Y(n_9783_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9784 (.A1(n_9557_o_0),
    .A2(n_9529_o_0),
    .B(n_9783_o_0),
    .C(n_9526_o_0),
    .Y(n_9784_o_0));
 AOI21xp33_ASAP7_75t_R n_9785 (.A1(n_9724_o_0),
    .A2(n_9636_o_0),
    .B(n_9417_o_0),
    .Y(n_9785_o_0));
 OAI31xp33_ASAP7_75t_R n_9786 (.A1(n_9508_o_0),
    .A2(n_9559_o_0),
    .A3(n_9643_o_0),
    .B(n_9785_o_0),
    .Y(n_9786_o_0));
 OAI21xp33_ASAP7_75t_R n_9787 (.A1(net85),
    .A2(n_9699_o_0),
    .B(n_9767_o_0),
    .Y(n_9787_o_0));
 NOR3xp33_ASAP7_75t_R n_9788 (.A(n_9787_o_0),
    .B(n_9619_o_0),
    .C(n_9542_o_0),
    .Y(n_9788_o_0));
 AOI321xp33_ASAP7_75t_R n_9789 (.A1(n_9716_o_0),
    .A2(n_9782_o_0),
    .A3(n_9633_o_0),
    .B1(n_9784_o_0),
    .B2(n_9786_o_0),
    .C(n_9788_o_0),
    .Y(n_9789_o_0));
 NAND2xp33_ASAP7_75t_R n_979 (.A(n_878_o_0),
    .B(n_882_o_0),
    .Y(n_979_o_0));
 INVx1_ASAP7_75t_R n_9790 (.A(n_9612_o_0),
    .Y(n_9790_o_0));
 NOR2xp33_ASAP7_75t_R n_9791 (.A(n_9609_o_0),
    .B(n_9613_o_0),
    .Y(n_9791_o_0));
 INVx1_ASAP7_75t_R n_9792 (.A(n_9783_o_0),
    .Y(n_9792_o_0));
 OAI21xp33_ASAP7_75t_R n_9793 (.A1(n_9558_o_0),
    .A2(n_9703_o_0),
    .B(n_9619_o_0),
    .Y(n_9793_o_0));
 OAI21xp33_ASAP7_75t_R n_9794 (.A1(n_9791_o_0),
    .A2(n_9792_o_0),
    .B(n_9793_o_0),
    .Y(n_9794_o_0));
 INVx1_ASAP7_75t_R n_9795 (.A(n_9563_o_0),
    .Y(n_9795_o_0));
 AOI31xp33_ASAP7_75t_R n_9796 (.A1(n_9558_o_0),
    .A2(n_9795_o_0),
    .A3(n_9531_o_0),
    .B(n_9417_o_0),
    .Y(n_9796_o_0));
 OAI21xp33_ASAP7_75t_R n_9797 (.A1(n_9616_o_0),
    .A2(n_9681_o_0),
    .B(n_9796_o_0),
    .Y(n_9797_o_0));
 AOI21xp33_ASAP7_75t_R n_9798 (.A1(n_9509_o_0),
    .A2(n_9762_o_0),
    .B(n_9619_o_0),
    .Y(n_9798_o_0));
 OAI31xp33_ASAP7_75t_R n_9799 (.A1(n_9574_o_0),
    .A2(n_9490_o_0),
    .A3(net85),
    .B(n_9798_o_0),
    .Y(n_9799_o_0));
 OAI21xp33_ASAP7_75t_R n_980 (.A1(key[18]),
    .A2(n_827_o_0),
    .B(n_834_o_0),
    .Y(n_980_o_0));
 AOI21xp33_ASAP7_75t_R n_9800 (.A1(n_9797_o_0),
    .A2(n_9799_o_0),
    .B(n_9542_o_0),
    .Y(n_9800_o_0));
 AOI311xp33_ASAP7_75t_R n_9801 (.A1(n_9542_o_0),
    .A2(n_9790_o_0),
    .A3(n_9794_o_0),
    .B(n_9721_o_0),
    .C(n_9800_o_0),
    .Y(n_9801_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9802 (.A1(n_9721_o_0),
    .A2(n_9789_o_0),
    .B(n_9801_o_0),
    .C(n_9544_o_0),
    .Y(n_9802_o_0));
 OAI21xp33_ASAP7_75t_R n_9803 (.A1(n_9422_o_0),
    .A2(n_9781_o_0),
    .B(n_9802_o_0),
    .Y(n_9803_o_0));
 INVx1_ASAP7_75t_R n_9804 (.A(n_9596_o_0),
    .Y(n_9804_o_0));
 NOR3xp33_ASAP7_75t_R n_9805 (.A(n_9652_o_0),
    .B(n_9616_o_0),
    .C(n_9508_o_0),
    .Y(n_9805_o_0));
 OAI21xp33_ASAP7_75t_R n_9806 (.A1(n_9575_o_0),
    .A2(n_9490_o_0),
    .B(n_9501_o_0),
    .Y(n_9806_o_0));
 OAI32xp33_ASAP7_75t_R n_9807 (.A1(n_9501_o_0),
    .A2(n_9804_o_0),
    .A3(n_9805_o_0),
    .B1(n_9806_o_0),
    .B2(n_9666_o_0),
    .Y(n_9807_o_0));
 AOI21xp33_ASAP7_75t_R n_9808 (.A1(n_9531_o_0),
    .A2(n_9595_o_0),
    .B(n_9558_o_0),
    .Y(n_9808_o_0));
 OAI21xp33_ASAP7_75t_R n_9809 (.A1(n_9531_o_0),
    .A2(n_9555_o_0),
    .B(n_9808_o_0),
    .Y(n_9809_o_0));
 INVx1_ASAP7_75t_R n_981 (.A(n_835_o_0),
    .Y(n_981_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9810 (.A1(n_9465_o_0),
    .A2(n_9603_o_0),
    .B(n_9655_o_0),
    .C(n_9542_o_0),
    .Y(n_9810_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9811 (.A1(n_9809_o_0),
    .A2(n_9571_o_0),
    .B(n_9542_o_0),
    .C(n_9810_o_0),
    .Y(n_9811_o_0));
 OAI21xp33_ASAP7_75t_R n_9812 (.A1(n_9544_o_0),
    .A2(n_9811_o_0),
    .B(n_9619_o_0),
    .Y(n_9812_o_0));
 AOI21xp33_ASAP7_75t_R n_9813 (.A1(n_9422_o_0),
    .A2(n_9807_o_0),
    .B(n_9812_o_0),
    .Y(n_9813_o_0));
 AOI211xp5_ASAP7_75t_R n_9814 (.A1(n_9604_o_0),
    .A2(n_9508_o_0),
    .B(n_9542_o_0),
    .C(n_9533_o_0),
    .Y(n_9814_o_0));
 NOR3xp33_ASAP7_75t_R n_9815 (.A(n_9616_o_0),
    .B(n_9529_o_0),
    .C(n_9508_o_0),
    .Y(n_9815_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9816 (.A1(n_9452_o_0),
    .A2(net26),
    .B(n_9577_o_0),
    .C(n_9558_o_0),
    .Y(n_9816_o_0));
 NOR3xp33_ASAP7_75t_R n_9817 (.A(n_9815_o_0),
    .B(n_9526_o_0),
    .C(n_9816_o_0),
    .Y(n_9817_o_0));
 INVx1_ASAP7_75t_R n_9818 (.A(n_9557_o_0),
    .Y(n_9818_o_0));
 OAI21xp33_ASAP7_75t_R n_9819 (.A1(n_9710_o_0),
    .A2(n_9699_o_0),
    .B(n_9523_o_0),
    .Y(n_9819_o_0));
 AOI211xp5_ASAP7_75t_R n_982 (.A1(n_980_o_0),
    .A2(n_981_o_0),
    .B(n_847_o_0),
    .C(n_864_o_0),
    .Y(n_982_o_0));
 OAI211xp5_ASAP7_75t_R n_9820 (.A1(n_9487_o_0),
    .A2(net2),
    .B(n_9488_o_0),
    .C(_00967_),
    .Y(n_9820_o_0));
 AOI22xp33_ASAP7_75t_R n_9821 (.A1(n_9531_o_0),
    .A2(n_9451_o_0),
    .B1(n_9820_o_0),
    .B2(n_9464_o_0),
    .Y(n_9821_o_0));
 AOI21xp33_ASAP7_75t_R n_9822 (.A1(n_9821_o_0),
    .A2(n_9509_o_0),
    .B(n_9542_o_0),
    .Y(n_9822_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9823 (.A1(n_9531_o_0),
    .A2(n_9508_o_0),
    .B(n_9822_o_0),
    .C(n_9422_o_0),
    .Y(n_9823_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9824 (.A1(n_9818_o_0),
    .A2(n_9564_o_0),
    .B(n_9819_o_0),
    .C(n_9823_o_0),
    .Y(n_9824_o_0));
 OAI31xp33_ASAP7_75t_R n_9825 (.A1(n_9660_o_0),
    .A2(n_9814_o_0),
    .A3(n_9817_o_0),
    .B(n_9824_o_0),
    .Y(n_9825_o_0));
 AO21x1_ASAP7_75t_R n_9826 (.A1(n_9825_o_0),
    .A2(n_9417_o_0),
    .B(n_9721_o_0),
    .Y(n_9826_o_0));
 OAI31xp33_ASAP7_75t_R n_9827 (.A1(n_9508_o_0),
    .A2(n_9555_o_0),
    .A3(n_9531_o_0),
    .B(n_9754_o_0),
    .Y(n_9827_o_0));
 INVx1_ASAP7_75t_R n_9828 (.A(n_9827_o_0),
    .Y(n_9828_o_0));
 NAND3xp33_ASAP7_75t_R n_9829 (.A(net22),
    .B(n_9465_o_0),
    .C(n_9435_o_0),
    .Y(n_9829_o_0));
 NAND2xp33_ASAP7_75t_R n_983 (.A(n_877_o_0),
    .B(n_982_o_0),
    .Y(n_983_o_0));
 NAND3xp33_ASAP7_75t_R n_9830 (.A(n_9828_o_0),
    .B(n_9829_o_0),
    .C(n_9523_o_0),
    .Y(n_9830_o_0));
 AOI21xp33_ASAP7_75t_R n_9831 (.A1(n_9531_o_0),
    .A2(n_9651_o_0),
    .B(n_9490_o_0),
    .Y(n_9831_o_0));
 AOI21xp33_ASAP7_75t_R n_9832 (.A1(n_9560_o_0),
    .A2(n_9831_o_0),
    .B(n_9542_o_0),
    .Y(n_9832_o_0));
 OAI21xp33_ASAP7_75t_R n_9833 (.A1(n_9615_o_0),
    .A2(n_9616_o_0),
    .B(n_9832_o_0),
    .Y(n_9833_o_0));
 NAND2xp33_ASAP7_75t_R n_9834 (.A(n_9435_o_0),
    .B(n_9591_o_0),
    .Y(n_9834_o_0));
 AOI22xp33_ASAP7_75t_R n_9835 (.A1(n_9647_o_0),
    .A2(n_9834_o_0),
    .B1(n_9680_o_0),
    .B2(n_9534_o_0),
    .Y(n_9835_o_0));
 OAI22xp33_ASAP7_75t_R n_9836 (.A1(n_9616_o_0),
    .A2(n_9508_o_0),
    .B1(n_9601_o_0),
    .B2(n_9435_o_0),
    .Y(n_9836_o_0));
 AOI21xp33_ASAP7_75t_R n_9837 (.A1(n_9542_o_0),
    .A2(n_9836_o_0),
    .B(n_9544_o_0),
    .Y(n_9837_o_0));
 OAI21xp33_ASAP7_75t_R n_9838 (.A1(n_9523_o_0),
    .A2(n_9835_o_0),
    .B(n_9837_o_0),
    .Y(n_9838_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9839 (.A1(n_9830_o_0),
    .A2(n_9833_o_0),
    .B(n_9567_o_0),
    .C(n_9838_o_0),
    .Y(n_9839_o_0));
 NOR2xp33_ASAP7_75t_R n_984 (.A(n_881_o_0),
    .B(n_935_o_0),
    .Y(n_984_o_0));
 OAI311xp33_ASAP7_75t_R n_9840 (.A1(net26),
    .A2(n_9435_o_0),
    .A3(n_9451_o_0),
    .B1(n_9671_o_0),
    .C1(n_9558_o_0),
    .Y(n_9840_o_0));
 OAI31xp33_ASAP7_75t_R n_9841 (.A1(n_9490_o_0),
    .A2(n_9510_o_0),
    .A3(n_9710_o_0),
    .B(n_9840_o_0),
    .Y(n_9841_o_0));
 INVx1_ASAP7_75t_R n_9842 (.A(n_9601_o_0),
    .Y(n_9842_o_0));
 AOI211xp5_ASAP7_75t_R n_9843 (.A1(n_9842_o_0),
    .A2(n_9531_o_0),
    .B(n_9699_o_0),
    .C(n_9523_o_0),
    .Y(n_9843_o_0));
 AO21x1_ASAP7_75t_R n_9844 (.A1(n_9542_o_0),
    .A2(n_9841_o_0),
    .B(n_9843_o_0),
    .Y(n_9844_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9845 (.A1(n_9588_o_0),
    .A2(n_9596_o_0),
    .B(n_9542_o_0),
    .C(n_9544_o_0),
    .Y(n_9845_o_0));
 NOR2xp33_ASAP7_75t_R n_9846 (.A(n_9609_o_0),
    .B(n_9602_o_0),
    .Y(n_9846_o_0));
 AO21x1_ASAP7_75t_R n_9847 (.A1(n_9846_o_0),
    .A2(n_9558_o_0),
    .B(n_9816_o_0),
    .Y(n_9847_o_0));
 INVx1_ASAP7_75t_R n_9848 (.A(n_9820_o_0),
    .Y(n_9848_o_0));
 OAI221xp5_ASAP7_75t_R n_9849 (.A1(n_9489_o_0),
    .A2(n_9848_o_0),
    .B1(n_9531_o_0),
    .B2(net26),
    .C(n_9532_o_0),
    .Y(n_9849_o_0));
 NAND2xp33_ASAP7_75t_R n_985 (.A(n_877_o_0),
    .B(n_984_o_0),
    .Y(n_985_o_0));
 OAI31xp33_ASAP7_75t_R n_9850 (.A1(n_9508_o_0),
    .A2(n_9528_o_0),
    .A3(n_9609_o_0),
    .B(n_9849_o_0),
    .Y(n_9850_o_0));
 AOI21xp33_ASAP7_75t_R n_9851 (.A1(n_9526_o_0),
    .A2(n_9850_o_0),
    .B(n_9544_o_0),
    .Y(n_9851_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9852 (.A1(n_9847_o_0),
    .A2(n_9501_o_0),
    .B(n_9851_o_0),
    .C(n_9416_o_1),
    .Y(n_9852_o_0));
 OAI21xp33_ASAP7_75t_R n_9853 (.A1(n_9844_o_0),
    .A2(n_9845_o_0),
    .B(n_9852_o_0),
    .Y(n_9853_o_0));
 OAI211xp5_ASAP7_75t_R n_9854 (.A1(n_9839_o_0),
    .A2(n_9632_o_0),
    .B(n_9853_o_0),
    .C(n_9600_o_0),
    .Y(n_9854_o_0));
 OA21x2_ASAP7_75t_R n_9855 (.A1(n_9813_o_0),
    .A2(n_9826_o_0),
    .B(n_9854_o_0),
    .Y(n_9855_o_0));
 NOR2xp33_ASAP7_75t_R n_9856 (.A(n_9452_o_0),
    .B(n_9508_o_0),
    .Y(n_9856_o_0));
 OA211x2_ASAP7_75t_R n_9857 (.A1(n_9530_o_0),
    .A2(n_9856_o_0),
    .B(n_9619_o_0),
    .C(n_9526_o_0),
    .Y(n_9857_o_0));
 OAI21xp33_ASAP7_75t_R n_9858 (.A1(n_9531_o_0),
    .A2(net22),
    .B(n_9680_o_0),
    .Y(n_9858_o_0));
 OAI31xp33_ASAP7_75t_R n_9859 (.A1(n_9508_o_0),
    .A2(n_9574_o_0),
    .A3(n_9569_o_0),
    .B(n_9858_o_0),
    .Y(n_9859_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_986 (.A1(n_979_o_0),
    .A2(n_983_o_0),
    .B(n_891_o_0),
    .C(n_985_o_0),
    .Y(n_986_o_0));
 OAI211xp5_ASAP7_75t_R n_9860 (.A1(n_9522_o_0),
    .A2(n_9521_o_0),
    .B(n_9859_o_0),
    .C(n_9417_o_0),
    .Y(n_9860_o_0));
 NAND3xp33_ASAP7_75t_R n_9861 (.A(n_9558_o_0),
    .B(n_9563_o_0),
    .C(n_9435_o_0),
    .Y(n_9861_o_0));
 OAI31xp33_ASAP7_75t_R n_9862 (.A1(n_9490_o_0),
    .A2(n_9569_o_0),
    .A3(n_9510_o_0),
    .B(n_9861_o_0),
    .Y(n_9862_o_0));
 NAND3xp33_ASAP7_75t_R n_9863 (.A(n_9862_o_0),
    .B(n_9542_o_0),
    .C(n_9417_o_0),
    .Y(n_9863_o_0));
 INVx1_ASAP7_75t_R n_9864 (.A(n_9416_o_0),
    .Y(n_9864_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9865 (.A1(net89),
    .A2(n_9519_o_0),
    .B(n_9435_o_0),
    .C(n_9682_o_0),
    .Y(n_9865_o_0));
 OAI31xp33_ASAP7_75t_R n_9866 (.A1(n_9490_o_0),
    .A2(n_9652_o_0),
    .A3(n_9616_o_0),
    .B(n_9865_o_0),
    .Y(n_9866_o_0));
 OAI211xp5_ASAP7_75t_R n_9867 (.A1(n_9864_o_0),
    .A2(n_9631_o_0),
    .B(n_9866_o_0),
    .C(n_9542_o_0),
    .Y(n_9867_o_0));
 NAND4xp25_ASAP7_75t_R n_9868 (.A(n_9860_o_0),
    .B(n_9863_o_0),
    .C(n_9867_o_0),
    .D(n_9660_o_0),
    .Y(n_9868_o_0));
 AOI22xp33_ASAP7_75t_R n_9869 (.A1(n_9570_o_0),
    .A2(n_9465_o_0),
    .B1(n_9558_o_0),
    .B2(n_9563_o_0),
    .Y(n_9869_o_0));
 INVx1_ASAP7_75t_R n_987 (.A(n_986_o_0),
    .Y(n_987_o_0));
 OAI311xp33_ASAP7_75t_R n_9870 (.A1(n_9435_o_0),
    .A2(n_9723_o_0),
    .A3(n_9722_o_0),
    .B1(n_9465_o_0),
    .C1(n_9509_o_0),
    .Y(n_9870_o_0));
 OAI31xp33_ASAP7_75t_R n_9871 (.A1(n_9508_o_0),
    .A2(n_9520_o_0),
    .A3(n_9607_o_0),
    .B(n_9870_o_0),
    .Y(n_9871_o_0));
 AOI21xp33_ASAP7_75t_R n_9872 (.A1(n_9542_o_0),
    .A2(n_9871_o_0),
    .B(n_9619_o_0),
    .Y(n_9872_o_0));
 OAI21xp33_ASAP7_75t_R n_9873 (.A1(n_9523_o_0),
    .A2(n_9869_o_0),
    .B(n_9872_o_0),
    .Y(n_9873_o_0));
 OA211x2_ASAP7_75t_R n_9874 (.A1(n_9508_o_0),
    .A2(n_9510_o_0),
    .B(n_9829_o_0),
    .C(n_9416_o_1),
    .Y(n_9874_o_0));
 AOI21xp33_ASAP7_75t_R n_9875 (.A1(n_9504_o_0),
    .A2(n_9570_o_0),
    .B(n_9762_o_0),
    .Y(n_9875_o_0));
 OAI22xp33_ASAP7_75t_R n_9876 (.A1(n_9874_o_0),
    .A2(n_9633_o_0),
    .B1(n_9523_o_0),
    .B2(n_9875_o_0),
    .Y(n_9876_o_0));
 AO21x1_ASAP7_75t_R n_9877 (.A1(n_9873_o_0),
    .A2(n_9876_o_0),
    .B(n_9567_o_0),
    .Y(n_9877_o_0));
 OAI21xp33_ASAP7_75t_R n_9878 (.A1(n_9857_o_0),
    .A2(n_9868_o_0),
    .B(n_9877_o_0),
    .Y(n_9878_o_0));
 OAI33xp33_ASAP7_75t_R n_9879 (.A1(n_9490_o_0),
    .A2(n_9602_o_0),
    .A3(n_9609_o_0),
    .B1(n_9555_o_0),
    .B2(n_9531_o_0),
    .B3(n_9508_o_0),
    .Y(n_9879_o_0));
 OAI211xp5_ASAP7_75t_R n_988 (.A1(net16),
    .A2(n_959_o_0),
    .B(n_987_o_0),
    .C(n_903_o_0),
    .Y(n_988_o_0));
 OAI21xp33_ASAP7_75t_R n_9880 (.A1(n_9435_o_0),
    .A2(n_9575_o_0),
    .B(n_9490_o_0),
    .Y(n_9880_o_0));
 OAI211xp5_ASAP7_75t_R n_9881 (.A1(n_9452_o_0),
    .A2(net26),
    .B(n_9453_o_0),
    .C(n_9465_o_0),
    .Y(n_9881_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9882 (.A1(n_9563_o_0),
    .A2(n_9435_o_0),
    .B(n_9880_o_0),
    .C(n_9881_o_0),
    .Y(n_9882_o_0));
 OAI21xp33_ASAP7_75t_R n_9883 (.A1(n_9417_o_0),
    .A2(n_9882_o_0),
    .B(n_9544_o_0),
    .Y(n_9883_o_0));
 INVx1_ASAP7_75t_R n_9884 (.A(n_9734_o_0),
    .Y(n_9884_o_0));
 AOI21xp33_ASAP7_75t_R n_9885 (.A1(n_9435_o_0),
    .A2(n_9563_o_0),
    .B(n_9558_o_0),
    .Y(n_9885_o_0));
 AOI22xp33_ASAP7_75t_R n_9886 (.A1(n_9696_o_0),
    .A2(n_9452_o_0),
    .B1(n_9884_o_0),
    .B2(n_9885_o_0),
    .Y(n_9886_o_0));
 NOR2xp33_ASAP7_75t_R n_9887 (.A(n_9531_o_0),
    .B(n_9483_o_0),
    .Y(n_9887_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9888 (.A1(n_9887_o_0),
    .A2(n_9808_o_0),
    .B(n_9632_o_0),
    .C(n_9422_o_0),
    .Y(n_9888_o_0));
 OAI21xp33_ASAP7_75t_R n_9889 (.A1(n_9417_o_0),
    .A2(n_9886_o_0),
    .B(n_9888_o_0),
    .Y(n_9889_o_0));
 NOR2xp33_ASAP7_75t_R n_989 (.A(n_859_o_0),
    .B(n_836_o_0),
    .Y(n_989_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9890 (.A1(n_9632_o_0),
    .A2(n_9879_o_0),
    .B(n_9883_o_0),
    .C(n_9889_o_0),
    .Y(n_9890_o_0));
 INVx1_ASAP7_75t_R n_9891 (.A(n_9890_o_0),
    .Y(n_9891_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9892 (.A1(n_9651_o_0),
    .A2(n_9435_o_0),
    .B(n_9491_o_0),
    .C(n_9572_o_0),
    .Y(n_9892_o_0));
 OA21x2_ASAP7_75t_R n_9893 (.A1(n_9753_o_0),
    .A2(n_9755_o_0),
    .B(n_9417_o_0),
    .Y(n_9893_o_0));
 AOI21xp33_ASAP7_75t_R n_9894 (.A1(n_9619_o_0),
    .A2(n_9892_o_0),
    .B(n_9893_o_0),
    .Y(n_9894_o_0));
 AOI211xp5_ASAP7_75t_R n_9895 (.A1(n_9558_o_0),
    .A2(net26),
    .B(n_9816_o_0),
    .C(n_9417_o_0),
    .Y(n_9895_o_0));
 OAI31xp33_ASAP7_75t_R n_9896 (.A1(n_9508_o_0),
    .A2(n_9520_o_0),
    .A3(n_9602_o_0),
    .B(n_9632_o_0),
    .Y(n_9896_o_0));
 OAI21xp33_ASAP7_75t_R n_9897 (.A1(n_9896_o_0),
    .A2(n_9700_o_0),
    .B(n_9544_o_0),
    .Y(n_9897_o_0));
 OAI21xp33_ASAP7_75t_R n_9898 (.A1(n_9895_o_0),
    .A2(n_9897_o_0),
    .B(n_9501_o_0),
    .Y(n_9898_o_0));
 AOI21xp33_ASAP7_75t_R n_9899 (.A1(n_9567_o_0),
    .A2(n_9894_o_0),
    .B(n_9898_o_0),
    .Y(n_9899_o_0));
 OAI211xp5_ASAP7_75t_R n_990 (.A1(n_847_o_0),
    .A2(n_859_o_0),
    .B(n_888_o_0),
    .C(n_836_o_0),
    .Y(n_990_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9900 (.A1(n_9891_o_0),
    .A2(n_9523_o_0),
    .B(n_9899_o_0),
    .C(n_9600_o_0),
    .Y(n_9900_o_0));
 OAI21xp33_ASAP7_75t_R n_9901 (.A1(n_9600_o_0),
    .A2(n_9878_o_0),
    .B(n_9900_o_0),
    .Y(n_9901_o_0));
 OAI21xp33_ASAP7_75t_R n_9902 (.A1(n_9435_o_0),
    .A2(n_9555_o_0),
    .B(n_9465_o_0),
    .Y(n_9902_o_0));
 NOR2xp33_ASAP7_75t_R n_9903 (.A(n_9602_o_0),
    .B(n_9902_o_0),
    .Y(n_9903_o_0));
 AOI31xp33_ASAP7_75t_R n_9904 (.A1(n_9558_o_0),
    .A2(n_9577_o_0),
    .A3(n_9492_o_0),
    .B(n_9903_o_0),
    .Y(n_9904_o_0));
 NAND2xp33_ASAP7_75t_R n_9905 (.A(n_9531_o_0),
    .B(n_9483_o_0),
    .Y(n_9905_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9906 (.A1(n_9595_o_0),
    .A2(n_9643_o_0),
    .B(n_9592_o_0),
    .C(n_9501_o_0),
    .Y(n_9906_o_0));
 AOI31xp33_ASAP7_75t_R n_9907 (.A1(n_9558_o_0),
    .A2(n_9905_o_0),
    .A3(n_9766_o_0),
    .B(n_9906_o_0),
    .Y(n_9907_o_0));
 OAI22xp33_ASAP7_75t_R n_9908 (.A1(n_9632_o_0),
    .A2(n_9904_o_0),
    .B1(n_9907_o_0),
    .B2(n_9633_o_0),
    .Y(n_9908_o_0));
 AOI21xp33_ASAP7_75t_R n_9909 (.A1(n_9558_o_0),
    .A2(n_9735_o_0),
    .B(n_9504_o_0),
    .Y(n_9909_o_0));
 NAND2xp33_ASAP7_75t_R n_991 (.A(n_877_o_0),
    .B(n_990_o_0),
    .Y(n_991_o_0));
 NAND3xp33_ASAP7_75t_R n_9910 (.A(n_9905_o_0),
    .B(n_9834_o_0),
    .C(n_9558_o_0),
    .Y(n_9910_o_0));
 OAI31xp33_ASAP7_75t_R n_9911 (.A1(n_9490_o_0),
    .A2(n_9795_o_0),
    .A3(n_9531_o_0),
    .B(n_9910_o_0),
    .Y(n_9911_o_0));
 AOI21xp33_ASAP7_75t_R n_9912 (.A1(n_9417_o_0),
    .A2(n_9911_o_0),
    .B(n_9526_o_0),
    .Y(n_9912_o_0));
 OAI21xp33_ASAP7_75t_R n_9913 (.A1(n_9909_o_0),
    .A2(n_9793_o_0),
    .B(n_9912_o_0),
    .Y(n_9913_o_0));
 OAI21xp33_ASAP7_75t_R n_9914 (.A1(n_9465_o_0),
    .A2(n_9538_o_0),
    .B(n_9542_o_0),
    .Y(n_9914_o_0));
 NOR2xp33_ASAP7_75t_R n_9915 (.A(n_9529_o_0),
    .B(n_9592_o_0),
    .Y(n_9915_o_0));
 NOR3xp33_ASAP7_75t_R n_9916 (.A(n_9508_o_0),
    .B(n_9531_o_0),
    .C(n_9451_o_0),
    .Y(n_9916_o_0));
 NOR2xp33_ASAP7_75t_R n_9917 (.A(n_9435_o_0),
    .B(n_9465_o_0),
    .Y(n_9917_o_0));
 AOI21xp33_ASAP7_75t_R n_9918 (.A1(n_9917_o_0),
    .A2(n_9842_o_0),
    .B(n_9523_o_0),
    .Y(n_9918_o_0));
 OAI321xp33_ASAP7_75t_R n_9919 (.A1(n_9531_o_0),
    .A2(n_9575_o_0),
    .A3(n_9508_o_0),
    .B1(n_9616_o_0),
    .B2(n_9663_o_0),
    .C(n_9918_o_0),
    .Y(n_9919_o_0));
 OA21x2_ASAP7_75t_R n_992 (.A1(n_989_o_0),
    .A2(n_877_o_0),
    .B(n_991_o_0),
    .Y(n_992_o_0));
 OAI31xp33_ASAP7_75t_R n_9920 (.A1(n_9914_o_0),
    .A2(n_9915_o_0),
    .A3(n_9916_o_0),
    .B(n_9919_o_0),
    .Y(n_9920_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9921 (.A1(n_9451_o_0),
    .A2(n_9591_o_0),
    .B(n_9652_o_0),
    .C(n_9490_o_0),
    .Y(n_9921_o_0));
 OAI21xp33_ASAP7_75t_R n_9922 (.A1(n_9591_o_0),
    .A2(n_9558_o_0),
    .B(n_9921_o_0),
    .Y(n_9922_o_0));
 OAI31xp33_ASAP7_75t_R n_9923 (.A1(n_9523_o_0),
    .A2(n_9922_o_0),
    .A3(n_9632_o_0),
    .B(n_9660_o_0),
    .Y(n_9923_o_0));
 NOR2xp33_ASAP7_75t_R n_9924 (.A(n_9531_o_0),
    .B(n_9508_o_0),
    .Y(n_9924_o_0));
 INVx1_ASAP7_75t_R n_9925 (.A(n_9746_o_0),
    .Y(n_9925_o_0));
 AOI211xp5_ASAP7_75t_R n_9926 (.A1(n_9842_o_0),
    .A2(n_9924_o_0),
    .B(n_9925_o_0),
    .C(n_9914_o_0),
    .Y(n_9926_o_0));
 AOI211xp5_ASAP7_75t_R n_9927 (.A1(n_9920_o_0),
    .A2(n_9417_o_0),
    .B(n_9923_o_0),
    .C(n_9926_o_0),
    .Y(n_9927_o_0));
 AOI31xp33_ASAP7_75t_R n_9928 (.A1(n_9544_o_0),
    .A2(n_9908_o_0),
    .A3(n_9913_o_0),
    .B(n_9927_o_0),
    .Y(n_9928_o_0));
 OAI21xp33_ASAP7_75t_R n_9929 (.A1(n_9531_o_0),
    .A2(net26),
    .B(n_9695_o_0),
    .Y(n_9929_o_0));
 NAND2xp33_ASAP7_75t_R n_993 (.A(n_836_o_0),
    .B(n_933_o_0),
    .Y(n_993_o_0));
 NOR3xp33_ASAP7_75t_R n_9930 (.A(n_9652_o_0),
    .B(n_9616_o_0),
    .C(n_9490_o_0),
    .Y(n_9930_o_0));
 AOI21xp33_ASAP7_75t_R n_9931 (.A1(n_9558_o_0),
    .A2(n_9929_o_0),
    .B(n_9930_o_0),
    .Y(n_9931_o_0));
 OAI21xp33_ASAP7_75t_R n_9932 (.A1(n_9452_o_0),
    .A2(n_9531_o_0),
    .B(n_9508_o_0),
    .Y(n_9932_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9933 (.A1(n_9531_o_0),
    .A2(n_9651_o_0),
    .B(n_9584_o_0),
    .C(n_9501_o_0),
    .Y(n_9933_o_0));
 AOI21xp33_ASAP7_75t_R n_9934 (.A1(n_9932_o_0),
    .A2(n_9933_o_0),
    .B(n_9417_o_0),
    .Y(n_9934_o_0));
 OAI31xp33_ASAP7_75t_R n_9935 (.A1(n_9508_o_0),
    .A2(n_9652_o_0),
    .A3(n_9616_o_0),
    .B(n_9613_o_0),
    .Y(n_9935_o_0));
 OAI21xp33_ASAP7_75t_R n_9936 (.A1(n_9522_o_0),
    .A2(n_9521_o_0),
    .B(n_9709_o_0),
    .Y(n_9936_o_0));
 OAI32xp33_ASAP7_75t_R n_9937 (.A1(n_9526_o_0),
    .A2(n_9619_o_0),
    .A3(n_9935_o_0),
    .B1(n_9936_o_0),
    .B2(n_9416_o_1),
    .Y(n_9937_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9938 (.A1(n_9523_o_0),
    .A2(n_9931_o_0),
    .B(n_9934_o_0),
    .C(n_9937_o_0),
    .Y(n_9938_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9939 (.A1(n_9558_o_0),
    .A2(n_9527_o_0),
    .B(n_9831_o_0),
    .C(n_9766_o_0),
    .Y(n_9939_o_0));
 INVx1_ASAP7_75t_R n_994 (.A(n_993_o_0),
    .Y(n_994_o_0));
 NAND3xp33_ASAP7_75t_R n_9940 (.A(n_9558_o_0),
    .B(n_9527_o_0),
    .C(n_9766_o_0),
    .Y(n_9940_o_0));
 OAI311xp33_ASAP7_75t_R n_9941 (.A1(n_9490_o_0),
    .A2(n_9652_o_0),
    .A3(n_9887_o_0),
    .B1(n_9501_o_0),
    .C1(n_9940_o_0),
    .Y(n_9941_o_0));
 OAI21xp33_ASAP7_75t_R n_9942 (.A1(n_9501_o_0),
    .A2(n_9939_o_0),
    .B(n_9941_o_0),
    .Y(n_9942_o_0));
 AOI22xp33_ASAP7_75t_R n_9943 (.A1(n_9504_o_0),
    .A2(n_9506_o_0),
    .B1(n_9558_o_0),
    .B2(n_9627_o_0),
    .Y(n_9943_o_0));
 OAI211xp5_ASAP7_75t_R n_9944 (.A1(n_9451_o_0),
    .A2(n_9531_o_0),
    .B(n_9754_o_0),
    .C(n_9490_o_0),
    .Y(n_9944_o_0));
 AOI31xp33_ASAP7_75t_R n_9945 (.A1(n_9501_o_0),
    .A2(n_9944_o_0),
    .A3(n_9902_o_0),
    .B(n_9619_o_0),
    .Y(n_9945_o_0));
 OAI21xp33_ASAP7_75t_R n_9946 (.A1(n_9501_o_0),
    .A2(n_9943_o_0),
    .B(n_9945_o_0),
    .Y(n_9946_o_0));
 OA211x2_ASAP7_75t_R n_9947 (.A1(n_9942_o_0),
    .A2(n_9417_o_0),
    .B(n_9567_o_0),
    .C(n_9946_o_0),
    .Y(n_9947_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9948 (.A1(n_9938_o_0),
    .A2(n_9544_o_0),
    .B(n_9947_o_0),
    .C(n_9553_o_0),
    .Y(n_9948_o_0));
 OAI21xp33_ASAP7_75t_R n_9949 (.A1(n_9661_o_0),
    .A2(n_9928_o_0),
    .B(n_9948_o_0),
    .Y(n_9949_o_0));
 OAI21xp33_ASAP7_75t_R n_995 (.A1(n_836_o_0),
    .A2(n_935_o_0),
    .B(n_877_o_0),
    .Y(n_995_o_0));
 OA21x2_ASAP7_75t_R n_9950 (.A1(n_9558_o_0),
    .A2(n_9595_o_0),
    .B(n_9921_o_0),
    .Y(n_9950_o_0));
 NAND2xp33_ASAP7_75t_R n_9951 (.A(n_9558_o_0),
    .B(n_9834_o_0),
    .Y(n_9951_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9952 (.A1(n_9490_o_0),
    .A2(n_9602_o_0),
    .B(n_9951_o_0),
    .C(n_9523_o_0),
    .Y(n_9952_o_0));
 AOI21xp33_ASAP7_75t_R n_9953 (.A1(n_9564_o_0),
    .A2(n_9952_o_0),
    .B(n_9619_o_0),
    .Y(n_9953_o_0));
 OAI21xp33_ASAP7_75t_R n_9954 (.A1(n_9501_o_0),
    .A2(n_9950_o_0),
    .B(n_9953_o_0),
    .Y(n_9954_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9955 (.A1(n_9531_o_0),
    .A2(n_9651_o_0),
    .B(n_9564_o_0),
    .C(n_9558_o_0),
    .Y(n_9955_o_0));
 OA21x2_ASAP7_75t_R n_9956 (.A1(n_9531_o_0),
    .A2(n_9795_o_0),
    .B(n_9584_o_0),
    .Y(n_9956_o_0));
 OAI21xp33_ASAP7_75t_R n_9957 (.A1(n_9955_o_0),
    .A2(n_9956_o_0),
    .B(n_9633_o_0),
    .Y(n_9957_o_0));
 NOR2xp33_ASAP7_75t_R n_9958 (.A(n_9531_o_0),
    .B(n_9651_o_0),
    .Y(n_9958_o_0));
 AOI211xp5_ASAP7_75t_R n_9959 (.A1(n_9762_o_0),
    .A2(n_9761_o_0),
    .B(n_9501_o_0),
    .C(n_9632_o_0),
    .Y(n_9959_o_0));
 NOR2xp33_ASAP7_75t_R n_996 (.A(n_836_o_0),
    .B(n_860_o_0),
    .Y(n_996_o_0));
 OAI31xp33_ASAP7_75t_R n_9960 (.A1(n_9490_o_0),
    .A2(n_9958_o_0),
    .A3(n_9609_o_0),
    .B(n_9959_o_0),
    .Y(n_9960_o_0));
 NAND4xp25_ASAP7_75t_R n_9961 (.A(n_9954_o_0),
    .B(n_9957_o_0),
    .C(n_9960_o_0),
    .D(n_9567_o_0),
    .Y(n_9961_o_0));
 OAI211xp5_ASAP7_75t_R n_9962 (.A1(n_9555_o_0),
    .A2(n_9435_o_0),
    .B(n_9560_o_0),
    .C(n_9558_o_0),
    .Y(n_9962_o_0));
 OAI31xp33_ASAP7_75t_R n_9963 (.A1(n_9574_o_0),
    .A2(n_9490_o_0),
    .A3(n_9652_o_0),
    .B(n_9962_o_0),
    .Y(n_9963_o_0));
 OAI21xp33_ASAP7_75t_R n_9964 (.A1(n_9508_o_0),
    .A2(n_9731_o_0),
    .B(n_9501_o_0),
    .Y(n_9964_o_0));
 NOR3xp33_ASAP7_75t_R n_9965 (.A(n_9559_o_0),
    .B(n_9539_o_0),
    .C(n_9490_o_0),
    .Y(n_9965_o_0));
 OAI21xp33_ASAP7_75t_R n_9966 (.A1(n_9964_o_0),
    .A2(n_9965_o_0),
    .B(n_9417_o_0),
    .Y(n_9966_o_0));
 NOR2xp33_ASAP7_75t_R n_9967 (.A(n_9508_o_0),
    .B(n_9575_o_0),
    .Y(n_9967_o_0));
 AOI211xp5_ASAP7_75t_R n_9968 (.A1(n_9587_o_0),
    .A2(n_9842_o_0),
    .B(n_9523_o_0),
    .C(n_9967_o_0),
    .Y(n_9968_o_0));
 AOI21xp33_ASAP7_75t_R n_9969 (.A1(n_9818_o_0),
    .A2(n_9905_o_0),
    .B(n_9819_o_0),
    .Y(n_9969_o_0));
 OAI21xp33_ASAP7_75t_R n_997 (.A1(n_994_o_0),
    .A2(n_996_o_0),
    .B(n_878_o_0),
    .Y(n_997_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9970 (.A1(n_9968_o_0),
    .A2(n_9969_o_0),
    .B(n_9416_o_1),
    .C(n_9660_o_0),
    .Y(n_9970_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9971 (.A1(n_9963_o_0),
    .A2(n_9542_o_0),
    .B(n_9966_o_0),
    .C(n_9970_o_0),
    .Y(n_9971_o_0));
 OA21x2_ASAP7_75t_R n_9972 (.A1(n_9435_o_0),
    .A2(n_9601_o_0),
    .B(n_9655_o_0),
    .Y(n_9972_o_0));
 AOI31xp33_ASAP7_75t_R n_9973 (.A1(n_9453_o_0),
    .A2(n_9465_o_0),
    .A3(n_9905_o_0),
    .B(n_9972_o_0),
    .Y(n_9973_o_0));
 OAI31xp33_ASAP7_75t_R n_9974 (.A1(n_9508_o_0),
    .A2(n_9576_o_0),
    .A3(n_9559_o_0),
    .B(n_9632_o_0),
    .Y(n_9974_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9975 (.A1(n_9453_o_0),
    .A2(n_9753_o_0),
    .B(n_9974_o_0),
    .C(n_9542_o_0),
    .Y(n_9975_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9976 (.A1(n_9616_o_0),
    .A2(n_9663_o_0),
    .B(n_9632_o_0),
    .C(n_9523_o_0),
    .Y(n_9976_o_0));
 NOR4xp25_ASAP7_75t_R n_9977 (.A(n_9699_o_0),
    .B(n_9505_o_0),
    .C(n_9523_o_0),
    .D(n_9416_o_1),
    .Y(n_9977_o_0));
 O2A1O1Ixp33_ASAP7_75t_R n_9978 (.A1(n_9831_o_0),
    .A2(n_9805_o_0),
    .B(n_9976_o_0),
    .C(n_9977_o_0),
    .Y(n_9978_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9979 (.A1(n_9973_o_0),
    .A2(n_9416_o_1),
    .B(n_9975_o_0),
    .C(n_9978_o_0),
    .Y(n_9979_o_0));
 OAI211xp5_ASAP7_75t_R n_998 (.A1(n_994_o_0),
    .A2(n_995_o_0),
    .B(n_997_o_0),
    .C(n_891_o_0),
    .Y(n_998_o_0));
 NAND3xp33_ASAP7_75t_R n_9980 (.A(n_9880_o_0),
    .B(n_9774_o_0),
    .C(n_9417_o_0),
    .Y(n_9980_o_0));
 OAI31xp33_ASAP7_75t_R n_9981 (.A1(n_9490_o_0),
    .A2(n_9958_o_0),
    .A3(n_9652_o_0),
    .B(n_9732_o_0),
    .Y(n_9981_o_0));
 AOI21xp33_ASAP7_75t_R n_9982 (.A1(n_9619_o_0),
    .A2(n_9981_o_0),
    .B(n_9542_o_0),
    .Y(n_9982_o_0));
 OAI21xp33_ASAP7_75t_R n_9983 (.A1(n_9902_o_0),
    .A2(n_9958_o_0),
    .B(n_9615_o_0),
    .Y(n_9983_o_0));
 OAI21xp33_ASAP7_75t_R n_9984 (.A1(n_9451_o_0),
    .A2(n_9558_o_0),
    .B(n_9619_o_0),
    .Y(n_9984_o_0));
 A2O1A1Ixp33_ASAP7_75t_R n_9985 (.A1(n_9834_o_0),
    .A2(n_9647_o_0),
    .B(n_9984_o_0),
    .C(n_9523_o_0),
    .Y(n_9985_o_0));
 AOI21xp33_ASAP7_75t_R n_9986 (.A1(n_9417_o_0),
    .A2(n_9983_o_0),
    .B(n_9985_o_0),
    .Y(n_9986_o_0));
 AOI21xp33_ASAP7_75t_R n_9987 (.A1(n_9980_o_0),
    .A2(n_9982_o_0),
    .B(n_9986_o_0),
    .Y(n_9987_o_0));
 OAI22xp33_ASAP7_75t_R n_9988 (.A1(n_9979_o_0),
    .A2(n_9544_o_0),
    .B1(n_9567_o_0),
    .B2(n_9987_o_0),
    .Y(n_9988_o_0));
 AOI32xp33_ASAP7_75t_R n_9989 (.A1(n_9961_o_0),
    .A2(n_9971_o_0),
    .A3(n_9600_o_0),
    .B1(n_9661_o_0),
    .B2(n_9988_o_0),
    .Y(n_9989_o_0));
 OAI21xp33_ASAP7_75t_R n_999 (.A1(net15),
    .A2(n_992_o_0),
    .B(n_998_o_0),
    .Y(n_999_o_0));
 INVx1_ASAP7_75t_R n_9990 (.A(_00866_),
    .Y(n_9990_o_0));
 XOR2xp5_ASAP7_75t_R n_9991 (.A(_01002_),
    .B(_01120_),
    .Y(n_9991_o_0));
 XNOR2xp5_ASAP7_75t_R n_9992 (.A(n_3136_o_0),
    .B(n_9991_o_0),
    .Y(n_9992_o_0));
 XNOR2xp5_ASAP7_75t_R n_9993 (.A(_01001_),
    .B(n_9992_o_0),
    .Y(n_9993_o_0));
 NAND2xp33_ASAP7_75t_R n_9994 (.A(_00665_),
    .B(net2),
    .Y(n_9994_o_0));
 OAI21xp33_ASAP7_75t_R n_9995 (.A1(net2),
    .A2(n_9993_o_0),
    .B(n_9994_o_0),
    .Y(n_9995_o_0));
 NOR2xp33_ASAP7_75t_R n_9996 (.A(n_9990_o_0),
    .B(n_9995_o_0),
    .Y(n_9996_o_0));
 AOI21xp33_ASAP7_75t_R n_9997 (.A1(n_9990_o_0),
    .A2(n_9995_o_0),
    .B(n_9996_o_0),
    .Y(n_9997_o_0));
 XNOR2xp5_ASAP7_75t_R n_9998 (.A(_01041_),
    .B(_01081_),
    .Y(n_9998_o_0));
 XNOR2xp5_ASAP7_75t_R n_9999 (.A(_01119_),
    .B(n_9998_o_0),
    .Y(n_9999_o_0));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_3247_o_0),
    .QN(_00996_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_3316_o_0),
    .QN(_00997_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_3367_o_0),
    .QN(_00998_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_3415_o_0),
    .QN(_00999_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_3457_o_0),
    .QN(_01000_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_3502_o_0),
    .QN(_01001_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_3552_o_0),
    .QN(_01002_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_3596_o_0),
    .QN(_01003_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_3831_o_0),
    .QN(_01004_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_3892_o_0),
    .QN(_01005_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_3952_o_0),
    .QN(_01006_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_4001_o_0),
    .QN(_01007_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_4052_o_0),
    .QN(_01008_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_4097_o_0),
    .QN(_01009_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_4143_o_0),
    .QN(_01010_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_4184_o_0),
    .QN(_01011_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_4444_o_0),
    .QN(_01012_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_4514_o_0),
    .QN(_01013_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_4574_o_0),
    .QN(_01014_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_4621_o_0),
    .QN(_01015_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_4668_o_0),
    .QN(_01016_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_4712_o_0),
    .QN(_01017_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_4758_o_0),
    .QN(_01018_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_4801_o_0),
    .QN(_01019_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_5096_o_0),
    .QN(_01020_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_5151_o_0),
    .QN(_01021_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_5215_o_0),
    .QN(_01022_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_5258_o_0),
    .QN(_01023_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_5299_o_0),
    .QN(_01024_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_5347_o_0),
    .QN(_01025_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_5394_o_0),
    .QN(_01026_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_5438_o_0),
    .QN(_01027_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_6189_o_0),
    .QN(_01036_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_6262_o_0),
    .QN(_01037_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_6320_o_0),
    .QN(_01038_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_6378_o_0),
    .QN(_01039_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_6425_o_0),
    .QN(_01040_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_6466_o_0),
    .QN(_01041_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_6508_o_0),
    .QN(_01042_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_6551_o_0),
    .QN(_01043_));
 DFFHQNx1_ASAP7_75t_R \sa10_sub[0]$_DFF_P_  (.CLK(clk),
    .D(n_5646_o_0),
    .QN(_01028_));
 DFFHQNx1_ASAP7_75t_R \sa10_sub[1]$_DFF_P_  (.CLK(clk),
    .D(n_5706_o_0),
    .QN(_01029_));
 DFFHQNx1_ASAP7_75t_R \sa10_sub[2]$_DFF_P_  (.CLK(clk),
    .D(n_5760_o_0),
    .QN(_01030_));
 DFFHQNx1_ASAP7_75t_R \sa10_sub[3]$_DFF_P_  (.CLK(clk),
    .D(n_5809_o_0),
    .QN(_01031_));
 DFFHQNx1_ASAP7_75t_R \sa10_sub[4]$_DFF_P_  (.CLK(clk),
    .D(n_5857_o_0),
    .QN(_01032_));
 DFFHQNx1_ASAP7_75t_R \sa10_sub[5]$_DFF_P_  (.CLK(clk),
    .D(n_5900_o_0),
    .QN(_01033_));
 DFFHQNx1_ASAP7_75t_R \sa10_sub[6]$_DFF_P_  (.CLK(clk),
    .D(n_5944_o_0),
    .QN(_01034_));
 DFFHQNx1_ASAP7_75t_R \sa10_sub[7]$_DFF_P_  (.CLK(clk),
    .D(n_5988_o_0),
    .QN(_01035_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_6755_o_0),
    .QN(_01044_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_6819_o_0),
    .QN(_01045_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_6887_o_0),
    .QN(_01046_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_6941_o_0),
    .QN(_01047_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_6985_o_0),
    .QN(_01048_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_7029_o_0),
    .QN(_01049_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_7072_o_0),
    .QN(_01050_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_7113_o_0),
    .QN(_01051_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_7330_o_0),
    .QN(_01052_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_7408_o_0),
    .QN(_01053_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_7468_o_0),
    .QN(_01054_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_7518_o_0),
    .QN(_01055_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_7563_o_0),
    .QN(_01056_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_7609_o_0),
    .QN(_01057_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_7655_o_0),
    .QN(_01058_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_7696_o_0),
    .QN(_01059_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_9069_o_0),
    .QN(_01076_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_9130_o_0),
    .QN(_01077_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_9190_o_0),
    .QN(_01078_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_9236_o_0),
    .QN(_01079_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_9281_o_0),
    .QN(_01080_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_9321_o_0),
    .QN(_01081_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_9369_o_0),
    .QN(_01082_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_9410_o_0),
    .QN(_00643_));
 DFFHQNx1_ASAP7_75t_R \sa20_sub[0]$_DFF_P_  (.CLK(clk),
    .D(n_7909_o_0),
    .QN(_01060_));
 DFFHQNx1_ASAP7_75t_R \sa20_sub[1]$_DFF_P_  (.CLK(clk),
    .D(n_7974_o_0),
    .QN(_01061_));
 DFFHQNx1_ASAP7_75t_R \sa20_sub[2]$_DFF_P_  (.CLK(clk),
    .D(n_8035_o_0),
    .QN(_01062_));
 DFFHQNx1_ASAP7_75t_R \sa20_sub[3]$_DFF_P_  (.CLK(clk),
    .D(n_8094_o_0),
    .QN(_01063_));
 DFFHQNx1_ASAP7_75t_R \sa20_sub[4]$_DFF_P_  (.CLK(clk),
    .D(n_8140_o_0),
    .QN(_01064_));
 DFFHQNx1_ASAP7_75t_R \sa20_sub[5]$_DFF_P_  (.CLK(clk),
    .D(n_8182_o_0),
    .QN(_01065_));
 DFFHQNx1_ASAP7_75t_R \sa20_sub[6]$_DFF_P_  (.CLK(clk),
    .D(n_8229_o_0),
    .QN(_01066_));
 DFFHQNx1_ASAP7_75t_R \sa20_sub[7]$_DFF_P_  (.CLK(clk),
    .D(n_8273_o_0),
    .QN(_01067_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_9623_o_0),
    .QN(_01083_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_9690_o_0),
    .QN(_01084_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_9752_o_0),
    .QN(_01085_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_9803_o_0),
    .QN(_01086_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_9855_o_0),
    .QN(_01087_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_9901_o_0),
    .QN(_01088_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_9949_o_0),
    .QN(_01089_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_9989_o_0),
    .QN(_01090_));
 DFFHQNx1_ASAP7_75t_R \sa21_sub[0]$_DFF_P_  (.CLK(clk),
    .D(n_8491_o_0),
    .QN(_01068_));
 DFFHQNx1_ASAP7_75t_R \sa21_sub[1]$_DFF_P_  (.CLK(clk),
    .D(n_8563_o_0),
    .QN(_01069_));
 DFFHQNx1_ASAP7_75t_R \sa21_sub[2]$_DFF_P_  (.CLK(clk),
    .D(n_8621_o_0),
    .QN(_01070_));
 DFFHQNx1_ASAP7_75t_R \sa21_sub[3]$_DFF_P_  (.CLK(clk),
    .D(n_8675_o_0),
    .QN(_01071_));
 DFFHQNx1_ASAP7_75t_R \sa21_sub[4]$_DFF_P_  (.CLK(clk),
    .D(n_8720_o_0),
    .QN(_01072_));
 DFFHQNx1_ASAP7_75t_R \sa21_sub[5]$_DFF_P_  (.CLK(clk),
    .D(n_8777_o_0),
    .QN(_01073_));
 DFFHQNx1_ASAP7_75t_R \sa21_sub[6]$_DFF_P_  (.CLK(clk),
    .D(n_8826_o_0),
    .QN(_01074_));
 DFFHQNx1_ASAP7_75t_R \sa21_sub[7]$_DFF_P_  (.CLK(clk),
    .D(n_8866_o_0),
    .QN(_01075_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[0]$_DFF_P_  (.CLK(clk),
    .D(n_11879_o_0),
    .QN(_01115_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[1]$_DFF_P_  (.CLK(clk),
    .D(n_11953_o_0),
    .QN(_01116_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[2]$_DFF_P_  (.CLK(clk),
    .D(n_12016_o_0),
    .QN(_01117_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[3]$_DFF_P_  (.CLK(clk),
    .D(n_12067_o_0),
    .QN(_01118_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[4]$_DFF_P_  (.CLK(clk),
    .D(n_12110_o_0),
    .QN(_01119_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[5]$_DFF_P_  (.CLK(clk),
    .D(n_12154_o_0),
    .QN(_01120_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[6]$_DFF_P_  (.CLK(clk),
    .D(n_12198_o_0),
    .QN(_01121_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[7]$_DFF_P_  (.CLK(clk),
    .D(n_12237_o_0),
    .QN(_00642_));
 DFFHQNx1_ASAP7_75t_R \sa30_sub[0]$_DFF_P_  (.CLK(clk),
    .D(n_10190_o_0),
    .QN(_01091_));
 DFFHQNx1_ASAP7_75t_R \sa30_sub[1]$_DFF_P_  (.CLK(clk),
    .D(n_10260_o_0),
    .QN(_01092_));
 DFFHQNx1_ASAP7_75t_R \sa30_sub[2]$_DFF_P_  (.CLK(clk),
    .D(n_10315_o_0),
    .QN(_01093_));
 DFFHQNx1_ASAP7_75t_R \sa30_sub[3]$_DFF_P_  (.CLK(clk),
    .D(n_10371_o_0),
    .QN(_01094_));
 DFFHQNx1_ASAP7_75t_R \sa30_sub[4]$_DFF_P_  (.CLK(clk),
    .D(n_10419_o_0),
    .QN(_01095_));
 DFFHQNx1_ASAP7_75t_R \sa30_sub[5]$_DFF_P_  (.CLK(clk),
    .D(n_10462_o_0),
    .QN(_01096_));
 DFFHQNx1_ASAP7_75t_R \sa30_sub[6]$_DFF_P_  (.CLK(clk),
    .D(n_10508_o_0),
    .QN(_01097_));
 DFFHQNx1_ASAP7_75t_R \sa30_sub[7]$_DFF_P_  (.CLK(clk),
    .D(n_10548_o_0),
    .QN(_01098_));
 DFFHQNx1_ASAP7_75t_R \sa31_sub[0]$_DFF_P_  (.CLK(clk),
    .D(n_10753_o_0),
    .QN(_01099_));
 DFFHQNx1_ASAP7_75t_R \sa31_sub[1]$_DFF_P_  (.CLK(clk),
    .D(n_10824_o_0),
    .QN(_01100_));
 DFFHQNx1_ASAP7_75t_R \sa31_sub[2]$_DFF_P_  (.CLK(clk),
    .D(n_10877_o_0),
    .QN(_01101_));
 DFFHQNx1_ASAP7_75t_R \sa31_sub[3]$_DFF_P_  (.CLK(clk),
    .D(n_10928_o_0),
    .QN(_01102_));
 DFFHQNx1_ASAP7_75t_R \sa31_sub[4]$_DFF_P_  (.CLK(clk),
    .D(n_10971_o_0),
    .QN(_01103_));
 DFFHQNx1_ASAP7_75t_R \sa31_sub[5]$_DFF_P_  (.CLK(clk),
    .D(n_11017_o_0),
    .QN(_01104_));
 DFFHQNx1_ASAP7_75t_R \sa31_sub[6]$_DFF_P_  (.CLK(clk),
    .D(n_11055_o_0),
    .QN(_01105_));
 DFFHQNx1_ASAP7_75t_R \sa31_sub[7]$_DFF_P_  (.CLK(clk),
    .D(n_11098_o_0),
    .QN(_01106_));
 DFFHQNx1_ASAP7_75t_R \sa32_sub[0]$_DFF_P_  (.CLK(clk),
    .D(n_11299_o_0),
    .QN(_01107_));
 DFFHQNx1_ASAP7_75t_R \sa32_sub[1]$_DFF_P_  (.CLK(clk),
    .D(n_11364_o_0),
    .QN(_01108_));
 DFFHQNx1_ASAP7_75t_R \sa32_sub[2]$_DFF_P_  (.CLK(clk),
    .D(n_11424_o_0),
    .QN(_01109_));
 DFFHQNx1_ASAP7_75t_R \sa32_sub[3]$_DFF_P_  (.CLK(clk),
    .D(n_11479_o_0),
    .QN(_01110_));
 DFFHQNx1_ASAP7_75t_R \sa32_sub[4]$_DFF_P_  (.CLK(clk),
    .D(n_11528_o_0),
    .QN(_01111_));
 DFFHQNx1_ASAP7_75t_R \sa32_sub[5]$_DFF_P_  (.CLK(clk),
    .D(n_11577_o_0),
    .QN(_01112_));
 DFFHQNx1_ASAP7_75t_R \sa32_sub[6]$_DFF_P_  (.CLK(clk),
    .D(n_11623_o_0),
    .QN(_01113_));
 DFFHQNx1_ASAP7_75t_R \sa32_sub[7]$_DFF_P_  (.CLK(clk),
    .D(n_11666_o_0),
    .QN(_01114_));
 BUFx6f_ASAP7_75t_R split (.A(_00858_),
    .Y(net));
 BUFx4f_ASAP7_75t_R split39 (.A(_00858_),
    .Y(net39));
 BUFx2_ASAP7_75t_R split49 (.A(n_11177_o_1),
    .Y(net49));
 BUFx2_ASAP7_75t_R split77 (.A(_00858_),
    .Y(net77));
 DFFHQNx1_ASAP7_75t_R \text_in_r[0]$_DFFE_PP_  (.CLK(clk),
    .D(n_12615_o_0),
    .QN(_00411_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[100]$_DFFE_PP_  (.CLK(clk),
    .D(n_12815_o_0),
    .QN(_00667_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[101]$_DFFE_PP_  (.CLK(clk),
    .D(n_12817_o_0),
    .QN(_00666_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[102]$_DFFE_PP_  (.CLK(clk),
    .D(n_12819_o_0),
    .QN(_00665_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[103]$_DFFE_PP_  (.CLK(clk),
    .D(n_12821_o_0),
    .QN(_00664_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[104]$_DFFE_PP_  (.CLK(clk),
    .D(n_12823_o_0),
    .QN(_00570_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[105]$_DFFE_PP_  (.CLK(clk),
    .D(n_12825_o_0),
    .QN(_00569_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[106]$_DFFE_PP_  (.CLK(clk),
    .D(n_12827_o_0),
    .QN(_00572_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[107]$_DFFE_PP_  (.CLK(clk),
    .D(n_12829_o_0),
    .QN(_00663_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[108]$_DFFE_PP_  (.CLK(clk),
    .D(n_12831_o_0),
    .QN(_00662_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[109]$_DFFE_PP_  (.CLK(clk),
    .D(n_12833_o_0),
    .QN(_00661_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[10]$_DFFE_PP_  (.CLK(clk),
    .D(n_12635_o_0),
    .QN(_00608_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[110]$_DFFE_PP_  (.CLK(clk),
    .D(n_12835_o_0),
    .QN(_00660_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[111]$_DFFE_PP_  (.CLK(clk),
    .D(n_12837_o_0),
    .QN(_00659_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[112]$_DFFE_PP_  (.CLK(clk),
    .D(n_12839_o_0),
    .QN(_00530_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[113]$_DFFE_PP_  (.CLK(clk),
    .D(n_12841_o_0),
    .QN(_00529_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[114]$_DFFE_PP_  (.CLK(clk),
    .D(n_12843_o_0),
    .QN(_00532_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[115]$_DFFE_PP_  (.CLK(clk),
    .D(n_12845_o_0),
    .QN(_00658_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[116]$_DFFE_PP_  (.CLK(clk),
    .D(n_12847_o_0),
    .QN(_00657_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[117]$_DFFE_PP_  (.CLK(clk),
    .D(n_12849_o_0),
    .QN(_00656_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[118]$_DFFE_PP_  (.CLK(clk),
    .D(n_12851_o_0),
    .QN(_00655_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[119]$_DFFE_PP_  (.CLK(clk),
    .D(n_12853_o_0),
    .QN(_00654_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[11]$_DFFE_PP_  (.CLK(clk),
    .D(n_12637_o_0),
    .QN(_00723_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[120]$_DFFE_PP_  (.CLK(clk),
    .D(n_12855_o_0),
    .QN(_00490_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[121]$_DFFE_PP_  (.CLK(clk),
    .D(n_12857_o_0),
    .QN(_00489_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[122]$_DFFE_PP_  (.CLK(clk),
    .D(n_12859_o_0),
    .QN(_00492_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[123]$_DFFE_PP_  (.CLK(clk),
    .D(n_12861_o_0),
    .QN(_00653_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[124]$_DFFE_PP_  (.CLK(clk),
    .D(n_12863_o_0),
    .QN(_00652_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[125]$_DFFE_PP_  (.CLK(clk),
    .D(n_12865_o_0),
    .QN(_00651_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[126]$_DFFE_PP_  (.CLK(clk),
    .D(n_12867_o_0),
    .QN(_00650_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[127]$_DFFE_PP_  (.CLK(clk),
    .D(n_12869_o_0),
    .QN(_00649_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[12]$_DFFE_PP_  (.CLK(clk),
    .D(n_12639_o_0),
    .QN(_00722_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[13]$_DFFE_PP_  (.CLK(clk),
    .D(n_12641_o_0),
    .QN(_00721_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[14]$_DFFE_PP_  (.CLK(clk),
    .D(n_12643_o_0),
    .QN(_00720_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[15]$_DFFE_PP_  (.CLK(clk),
    .D(n_12645_o_0),
    .QN(_00719_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[16]$_DFFE_PP_  (.CLK(clk),
    .D(n_12647_o_0),
    .QN(_00560_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[17]$_DFFE_PP_  (.CLK(clk),
    .D(n_12649_o_0),
    .QN(_00559_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[18]$_DFFE_PP_  (.CLK(clk),
    .D(n_12651_o_0),
    .QN(_00562_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[19]$_DFFE_PP_  (.CLK(clk),
    .D(n_12653_o_0),
    .QN(_00718_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[1]$_DFFE_PP_  (.CLK(clk),
    .D(n_12617_o_0),
    .QN(_00410_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[20]$_DFFE_PP_  (.CLK(clk),
    .D(n_12655_o_0),
    .QN(_00717_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[21]$_DFFE_PP_  (.CLK(clk),
    .D(n_12657_o_0),
    .QN(_00716_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[22]$_DFFE_PP_  (.CLK(clk),
    .D(n_12659_o_0),
    .QN(_00715_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[23]$_DFFE_PP_  (.CLK(clk),
    .D(n_12661_o_0),
    .QN(_00714_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[24]$_DFFE_PP_  (.CLK(clk),
    .D(n_12663_o_0),
    .QN(_00520_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[25]$_DFFE_PP_  (.CLK(clk),
    .D(n_12665_o_0),
    .QN(_00519_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[26]$_DFFE_PP_  (.CLK(clk),
    .D(n_12667_o_0),
    .QN(_00522_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[27]$_DFFE_PP_  (.CLK(clk),
    .D(n_12669_o_0),
    .QN(_00713_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[28]$_DFFE_PP_  (.CLK(clk),
    .D(n_12671_o_0),
    .QN(_00712_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[29]$_DFFE_PP_  (.CLK(clk),
    .D(n_12673_o_0),
    .QN(_00711_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[2]$_DFFE_PP_  (.CLK(clk),
    .D(n_12619_o_0),
    .QN(_00413_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[30]$_DFFE_PP_  (.CLK(clk),
    .D(n_12675_o_0),
    .QN(_00710_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[31]$_DFFE_PP_  (.CLK(clk),
    .D(n_12677_o_0),
    .QN(_00709_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[32]$_DFFE_PP_  (.CLK(clk),
    .D(n_12679_o_0),
    .QN(_00638_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[33]$_DFFE_PP_  (.CLK(clk),
    .D(n_12681_o_0),
    .QN(_00637_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[34]$_DFFE_PP_  (.CLK(clk),
    .D(n_12683_o_0),
    .QN(_00639_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[35]$_DFFE_PP_  (.CLK(clk),
    .D(n_12685_o_0),
    .QN(_00708_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[36]$_DFFE_PP_  (.CLK(clk),
    .D(n_12687_o_0),
    .QN(_00707_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[37]$_DFFE_PP_  (.CLK(clk),
    .D(n_12689_o_0),
    .QN(_00706_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[38]$_DFFE_PP_  (.CLK(clk),
    .D(n_12691_o_0),
    .QN(_00705_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[39]$_DFFE_PP_  (.CLK(clk),
    .D(n_12693_o_0),
    .QN(_00704_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[3]$_DFFE_PP_  (.CLK(clk),
    .D(n_12621_o_0),
    .QN(_00728_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[40]$_DFFE_PP_  (.CLK(clk),
    .D(n_12695_o_0),
    .QN(_00594_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[41]$_DFFE_PP_  (.CLK(clk),
    .D(n_12697_o_0),
    .QN(_00593_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[42]$_DFFE_PP_  (.CLK(clk),
    .D(n_12699_o_0),
    .QN(_00596_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[43]$_DFFE_PP_  (.CLK(clk),
    .D(n_12701_o_0),
    .QN(_00703_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[44]$_DFFE_PP_  (.CLK(clk),
    .D(n_12703_o_0),
    .QN(_00702_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[45]$_DFFE_PP_  (.CLK(clk),
    .D(n_12705_o_0),
    .QN(_00701_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[46]$_DFFE_PP_  (.CLK(clk),
    .D(n_12707_o_0),
    .QN(_00700_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[47]$_DFFE_PP_  (.CLK(clk),
    .D(n_12709_o_0),
    .QN(_00699_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[48]$_DFFE_PP_  (.CLK(clk),
    .D(n_12711_o_0),
    .QN(_00550_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[49]$_DFFE_PP_  (.CLK(clk),
    .D(n_12713_o_0),
    .QN(_00549_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[4]$_DFFE_PP_  (.CLK(clk),
    .D(n_12623_o_0),
    .QN(_00727_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[50]$_DFFE_PP_  (.CLK(clk),
    .D(n_12715_o_0),
    .QN(_00552_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[51]$_DFFE_PP_  (.CLK(clk),
    .D(n_12717_o_0),
    .QN(_00698_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[52]$_DFFE_PP_  (.CLK(clk),
    .D(n_12719_o_0),
    .QN(_00697_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[53]$_DFFE_PP_  (.CLK(clk),
    .D(n_12721_o_0),
    .QN(_00696_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[54]$_DFFE_PP_  (.CLK(clk),
    .D(n_12723_o_0),
    .QN(_00695_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[55]$_DFFE_PP_  (.CLK(clk),
    .D(n_12725_o_0),
    .QN(_00694_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[56]$_DFFE_PP_  (.CLK(clk),
    .D(n_12727_o_0),
    .QN(_00510_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[57]$_DFFE_PP_  (.CLK(clk),
    .D(n_12729_o_0),
    .QN(_00509_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[58]$_DFFE_PP_  (.CLK(clk),
    .D(n_12731_o_0),
    .QN(_00512_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[59]$_DFFE_PP_  (.CLK(clk),
    .D(n_12733_o_0),
    .QN(_00693_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[5]$_DFFE_PP_  (.CLK(clk),
    .D(n_12625_o_0),
    .QN(_00726_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[60]$_DFFE_PP_  (.CLK(clk),
    .D(n_12735_o_0),
    .QN(_00692_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[61]$_DFFE_PP_  (.CLK(clk),
    .D(n_12737_o_0),
    .QN(_00691_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[62]$_DFFE_PP_  (.CLK(clk),
    .D(n_12739_o_0),
    .QN(_00690_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[63]$_DFFE_PP_  (.CLK(clk),
    .D(n_12741_o_0),
    .QN(_00689_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[64]$_DFFE_PP_  (.CLK(clk),
    .D(n_12743_o_0),
    .QN(_00628_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[65]$_DFFE_PP_  (.CLK(clk),
    .D(n_12745_o_0),
    .QN(_00627_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[66]$_DFFE_PP_  (.CLK(clk),
    .D(n_12747_o_0),
    .QN(_00630_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[67]$_DFFE_PP_  (.CLK(clk),
    .D(n_12749_o_0),
    .QN(_00688_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[68]$_DFFE_PP_  (.CLK(clk),
    .D(n_12751_o_0),
    .QN(_00687_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[69]$_DFFE_PP_  (.CLK(clk),
    .D(n_12753_o_0),
    .QN(_00686_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[6]$_DFFE_PP_  (.CLK(clk),
    .D(n_12627_o_0),
    .QN(_00725_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[70]$_DFFE_PP_  (.CLK(clk),
    .D(n_12755_o_0),
    .QN(_00685_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[71]$_DFFE_PP_  (.CLK(clk),
    .D(n_12757_o_0),
    .QN(_00684_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[72]$_DFFE_PP_  (.CLK(clk),
    .D(n_12759_o_0),
    .QN(_00582_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[73]$_DFFE_PP_  (.CLK(clk),
    .D(n_12761_o_0),
    .QN(_00581_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[74]$_DFFE_PP_  (.CLK(clk),
    .D(n_12763_o_0),
    .QN(_00584_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[75]$_DFFE_PP_  (.CLK(clk),
    .D(n_12765_o_0),
    .QN(_00683_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[76]$_DFFE_PP_  (.CLK(clk),
    .D(n_12767_o_0),
    .QN(_00682_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[77]$_DFFE_PP_  (.CLK(clk),
    .D(n_12769_o_0),
    .QN(_00681_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[78]$_DFFE_PP_  (.CLK(clk),
    .D(n_12771_o_0),
    .QN(_00680_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[79]$_DFFE_PP_  (.CLK(clk),
    .D(n_12773_o_0),
    .QN(_00679_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[7]$_DFFE_PP_  (.CLK(clk),
    .D(n_12629_o_0),
    .QN(_00724_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[80]$_DFFE_PP_  (.CLK(clk),
    .D(n_12775_o_0),
    .QN(_00540_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[81]$_DFFE_PP_  (.CLK(clk),
    .D(n_12777_o_0),
    .QN(_00539_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[82]$_DFFE_PP_  (.CLK(clk),
    .D(n_12779_o_0),
    .QN(_00542_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[83]$_DFFE_PP_  (.CLK(clk),
    .D(n_12781_o_0),
    .QN(_00678_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[84]$_DFFE_PP_  (.CLK(clk),
    .D(n_12783_o_0),
    .QN(_00677_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[85]$_DFFE_PP_  (.CLK(clk),
    .D(n_12785_o_0),
    .QN(_00676_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[86]$_DFFE_PP_  (.CLK(clk),
    .D(n_12787_o_0),
    .QN(_00675_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[87]$_DFFE_PP_  (.CLK(clk),
    .D(n_12789_o_0),
    .QN(_00674_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[88]$_DFFE_PP_  (.CLK(clk),
    .D(n_12791_o_0),
    .QN(_00500_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[89]$_DFFE_PP_  (.CLK(clk),
    .D(n_12793_o_0),
    .QN(_00499_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[8]$_DFFE_PP_  (.CLK(clk),
    .D(n_12631_o_0),
    .QN(_00606_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[90]$_DFFE_PP_  (.CLK(clk),
    .D(n_12795_o_0),
    .QN(_00502_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[91]$_DFFE_PP_  (.CLK(clk),
    .D(n_12797_o_0),
    .QN(_00673_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[92]$_DFFE_PP_  (.CLK(clk),
    .D(n_12799_o_0),
    .QN(_00672_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[93]$_DFFE_PP_  (.CLK(clk),
    .D(n_12801_o_0),
    .QN(_00671_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[94]$_DFFE_PP_  (.CLK(clk),
    .D(n_12803_o_0),
    .QN(_00670_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[95]$_DFFE_PP_  (.CLK(clk),
    .D(n_12805_o_0),
    .QN(_00669_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[96]$_DFFE_PP_  (.CLK(clk),
    .D(n_12807_o_0),
    .QN(_00618_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[97]$_DFFE_PP_  (.CLK(clk),
    .D(n_12809_o_0),
    .QN(_00617_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[98]$_DFFE_PP_  (.CLK(clk),
    .D(n_12811_o_0),
    .QN(_00620_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[99]$_DFFE_PP_  (.CLK(clk),
    .D(n_12813_o_0),
    .QN(_00668_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[9]$_DFFE_PP_  (.CLK(clk),
    .D(n_12633_o_0),
    .QN(_00605_));
 DFFHQNx1_ASAP7_75t_R \text_out[0]$_DFF_P_  (.CLK(clk),
    .D(n_12346_o_0),
    .QN(_00730_));
 DFFHQNx1_ASAP7_75t_R \text_out[100]$_DFF_P_  (.CLK(clk),
    .D(n_12246_o_0),
    .QN(_00758_));
 DFFHQNx1_ASAP7_75t_R \text_out[101]$_DFF_P_  (.CLK(clk),
    .D(n_12247_o_0),
    .QN(_00759_));
 DFFHQNx1_ASAP7_75t_R \text_out[102]$_DFF_P_  (.CLK(clk),
    .D(n_12248_o_0),
    .QN(_00760_));
 DFFHQNx1_ASAP7_75t_R \text_out[103]$_DFF_P_  (.CLK(clk),
    .D(n_12249_o_0),
    .QN(_00761_));
 DFFHQNx1_ASAP7_75t_R \text_out[104]$_DFF_P_  (.CLK(clk),
    .D(n_12250_o_0),
    .QN(_00786_));
 DFFHQNx1_ASAP7_75t_R \text_out[105]$_DFF_P_  (.CLK(clk),
    .D(n_12251_o_0),
    .QN(_00787_));
 DFFHQNx1_ASAP7_75t_R \text_out[106]$_DFF_P_  (.CLK(clk),
    .D(n_12252_o_0),
    .QN(_00788_));
 DFFHQNx1_ASAP7_75t_R \text_out[107]$_DFF_P_  (.CLK(clk),
    .D(n_12253_o_0),
    .QN(_00789_));
 DFFHQNx1_ASAP7_75t_R \text_out[108]$_DFF_P_  (.CLK(clk),
    .D(n_12254_o_0),
    .QN(_00790_));
 DFFHQNx1_ASAP7_75t_R \text_out[109]$_DFF_P_  (.CLK(clk),
    .D(n_12255_o_0),
    .QN(_00791_));
 DFFHQNx1_ASAP7_75t_R \text_out[10]$_DFF_P_  (.CLK(clk),
    .D(n_12276_o_0),
    .QN(_00764_));
 DFFHQNx1_ASAP7_75t_R \text_out[110]$_DFF_P_  (.CLK(clk),
    .D(n_12256_o_0),
    .QN(_00792_));
 DFFHQNx1_ASAP7_75t_R \text_out[111]$_DFF_P_  (.CLK(clk),
    .D(n_12257_o_0),
    .QN(_00793_));
 DFFHQNx1_ASAP7_75t_R \text_out[112]$_DFF_P_  (.CLK(clk),
    .D(n_12258_o_0),
    .QN(_00818_));
 DFFHQNx1_ASAP7_75t_R \text_out[113]$_DFF_P_  (.CLK(clk),
    .D(n_12259_o_0),
    .QN(_00819_));
 DFFHQNx1_ASAP7_75t_R \text_out[114]$_DFF_P_  (.CLK(clk),
    .D(n_12260_o_0),
    .QN(_00820_));
 DFFHQNx1_ASAP7_75t_R \text_out[115]$_DFF_P_  (.CLK(clk),
    .D(n_12261_o_0),
    .QN(_00821_));
 DFFHQNx1_ASAP7_75t_R \text_out[116]$_DFF_P_  (.CLK(clk),
    .D(n_12262_o_0),
    .QN(_00822_));
 DFFHQNx1_ASAP7_75t_R \text_out[117]$_DFF_P_  (.CLK(clk),
    .D(n_12263_o_0),
    .QN(_00823_));
 DFFHQNx1_ASAP7_75t_R \text_out[118]$_DFF_P_  (.CLK(clk),
    .D(n_12264_o_0),
    .QN(_00824_));
 DFFHQNx1_ASAP7_75t_R \text_out[119]$_DFF_P_  (.CLK(clk),
    .D(n_12265_o_0),
    .QN(_00825_));
 DFFHQNx1_ASAP7_75t_R \text_out[11]$_DFF_P_  (.CLK(clk),
    .D(n_12277_o_0),
    .QN(_00765_));
 DFFHQNx1_ASAP7_75t_R \text_out[120]$_DFF_P_  (.CLK(clk),
    .D(n_12266_o_0),
    .QN(_00850_));
 DFFHQNx1_ASAP7_75t_R \text_out[121]$_DFF_P_  (.CLK(clk),
    .D(n_12267_o_0),
    .QN(_00851_));
 DFFHQNx1_ASAP7_75t_R \text_out[122]$_DFF_P_  (.CLK(clk),
    .D(n_12268_o_0),
    .QN(_00852_));
 DFFHQNx1_ASAP7_75t_R \text_out[123]$_DFF_P_  (.CLK(clk),
    .D(n_12269_o_0),
    .QN(_00853_));
 DFFHQNx1_ASAP7_75t_R \text_out[124]$_DFF_P_  (.CLK(clk),
    .D(n_12270_o_0),
    .QN(_00854_));
 DFFHQNx1_ASAP7_75t_R \text_out[125]$_DFF_P_  (.CLK(clk),
    .D(n_12271_o_0),
    .QN(_00855_));
 DFFHQNx1_ASAP7_75t_R \text_out[126]$_DFF_P_  (.CLK(clk),
    .D(n_12272_o_0),
    .QN(_00856_));
 DFFHQNx1_ASAP7_75t_R \text_out[127]$_DFF_P_  (.CLK(clk),
    .D(n_12273_o_0),
    .QN(_00857_));
 DFFHQNx1_ASAP7_75t_R \text_out[12]$_DFF_P_  (.CLK(clk),
    .D(n_12278_o_0),
    .QN(_00766_));
 DFFHQNx1_ASAP7_75t_R \text_out[13]$_DFF_P_  (.CLK(clk),
    .D(n_12279_o_0),
    .QN(_00767_));
 DFFHQNx1_ASAP7_75t_R \text_out[14]$_DFF_P_  (.CLK(clk),
    .D(n_12280_o_0),
    .QN(_00768_));
 DFFHQNx1_ASAP7_75t_R \text_out[15]$_DFF_P_  (.CLK(clk),
    .D(n_12281_o_0),
    .QN(_00769_));
 DFFHQNx1_ASAP7_75t_R \text_out[16]$_DFF_P_  (.CLK(clk),
    .D(n_12282_o_0),
    .QN(_00794_));
 DFFHQNx1_ASAP7_75t_R \text_out[17]$_DFF_P_  (.CLK(clk),
    .D(n_12283_o_0),
    .QN(_00795_));
 DFFHQNx1_ASAP7_75t_R \text_out[18]$_DFF_P_  (.CLK(clk),
    .D(n_12284_o_0),
    .QN(_00796_));
 DFFHQNx1_ASAP7_75t_R \text_out[19]$_DFF_P_  (.CLK(clk),
    .D(n_12285_o_0),
    .QN(_00797_));
 DFFHQNx1_ASAP7_75t_R \text_out[1]$_DFF_P_  (.CLK(clk),
    .D(n_12347_o_0),
    .QN(_00731_));
 DFFHQNx1_ASAP7_75t_R \text_out[20]$_DFF_P_  (.CLK(clk),
    .D(n_12286_o_0),
    .QN(_00798_));
 DFFHQNx1_ASAP7_75t_R \text_out[21]$_DFF_P_  (.CLK(clk),
    .D(n_12287_o_0),
    .QN(_00799_));
 DFFHQNx1_ASAP7_75t_R \text_out[22]$_DFF_P_  (.CLK(clk),
    .D(n_12288_o_0),
    .QN(_00800_));
 DFFHQNx1_ASAP7_75t_R \text_out[23]$_DFF_P_  (.CLK(clk),
    .D(n_12289_o_0),
    .QN(_00801_));
 DFFHQNx1_ASAP7_75t_R \text_out[24]$_DFF_P_  (.CLK(clk),
    .D(n_12290_o_0),
    .QN(_00826_));
 DFFHQNx1_ASAP7_75t_R \text_out[25]$_DFF_P_  (.CLK(clk),
    .D(n_12291_o_0),
    .QN(_00827_));
 DFFHQNx1_ASAP7_75t_R \text_out[26]$_DFF_P_  (.CLK(clk),
    .D(n_12292_o_0),
    .QN(_00828_));
 DFFHQNx1_ASAP7_75t_R \text_out[27]$_DFF_P_  (.CLK(clk),
    .D(n_12293_o_0),
    .QN(_00829_));
 DFFHQNx1_ASAP7_75t_R \text_out[28]$_DFF_P_  (.CLK(clk),
    .D(n_12294_o_0),
    .QN(_00830_));
 DFFHQNx1_ASAP7_75t_R \text_out[29]$_DFF_P_  (.CLK(clk),
    .D(n_12295_o_0),
    .QN(_00831_));
 DFFHQNx1_ASAP7_75t_R \text_out[2]$_DFF_P_  (.CLK(clk),
    .D(n_12348_o_0),
    .QN(_00732_));
 DFFHQNx1_ASAP7_75t_R \text_out[30]$_DFF_P_  (.CLK(clk),
    .D(n_12296_o_0),
    .QN(_00832_));
 DFFHQNx1_ASAP7_75t_R \text_out[31]$_DFF_P_  (.CLK(clk),
    .D(n_12297_o_0),
    .QN(_00833_));
 DFFHQNx1_ASAP7_75t_R \text_out[32]$_DFF_P_  (.CLK(clk),
    .D(n_12298_o_0),
    .QN(_00738_));
 DFFHQNx1_ASAP7_75t_R \text_out[33]$_DFF_P_  (.CLK(clk),
    .D(n_12299_o_0),
    .QN(_00739_));
 DFFHQNx1_ASAP7_75t_R \text_out[34]$_DFF_P_  (.CLK(clk),
    .D(n_12300_o_0),
    .QN(_00740_));
 DFFHQNx1_ASAP7_75t_R \text_out[35]$_DFF_P_  (.CLK(clk),
    .D(n_12301_o_0),
    .QN(_00741_));
 DFFHQNx1_ASAP7_75t_R \text_out[36]$_DFF_P_  (.CLK(clk),
    .D(n_12302_o_0),
    .QN(_00742_));
 DFFHQNx1_ASAP7_75t_R \text_out[37]$_DFF_P_  (.CLK(clk),
    .D(n_12303_o_0),
    .QN(_00743_));
 DFFHQNx1_ASAP7_75t_R \text_out[38]$_DFF_P_  (.CLK(clk),
    .D(n_12304_o_0),
    .QN(_00744_));
 DFFHQNx1_ASAP7_75t_R \text_out[39]$_DFF_P_  (.CLK(clk),
    .D(n_12305_o_0),
    .QN(_00745_));
 DFFHQNx1_ASAP7_75t_R \text_out[3]$_DFF_P_  (.CLK(clk),
    .D(n_12349_o_0),
    .QN(_00733_));
 DFFHQNx1_ASAP7_75t_R \text_out[40]$_DFF_P_  (.CLK(clk),
    .D(n_12306_o_0),
    .QN(_00770_));
 DFFHQNx1_ASAP7_75t_R \text_out[41]$_DFF_P_  (.CLK(clk),
    .D(n_12307_o_0),
    .QN(_00771_));
 DFFHQNx1_ASAP7_75t_R \text_out[42]$_DFF_P_  (.CLK(clk),
    .D(n_12308_o_0),
    .QN(_00772_));
 DFFHQNx1_ASAP7_75t_R \text_out[43]$_DFF_P_  (.CLK(clk),
    .D(n_12309_o_0),
    .QN(_00773_));
 DFFHQNx1_ASAP7_75t_R \text_out[44]$_DFF_P_  (.CLK(clk),
    .D(n_12310_o_0),
    .QN(_00774_));
 DFFHQNx1_ASAP7_75t_R \text_out[45]$_DFF_P_  (.CLK(clk),
    .D(n_12311_o_0),
    .QN(_00775_));
 DFFHQNx1_ASAP7_75t_R \text_out[46]$_DFF_P_  (.CLK(clk),
    .D(n_12312_o_0),
    .QN(_00776_));
 DFFHQNx1_ASAP7_75t_R \text_out[47]$_DFF_P_  (.CLK(clk),
    .D(n_12313_o_0),
    .QN(_00777_));
 DFFHQNx1_ASAP7_75t_R \text_out[48]$_DFF_P_  (.CLK(clk),
    .D(n_12314_o_0),
    .QN(_00802_));
 DFFHQNx1_ASAP7_75t_R \text_out[49]$_DFF_P_  (.CLK(clk),
    .D(n_12315_o_0),
    .QN(_00803_));
 DFFHQNx1_ASAP7_75t_R \text_out[4]$_DFF_P_  (.CLK(clk),
    .D(n_12350_o_0),
    .QN(_00734_));
 DFFHQNx1_ASAP7_75t_R \text_out[50]$_DFF_P_  (.CLK(clk),
    .D(n_12316_o_0),
    .QN(_00804_));
 DFFHQNx1_ASAP7_75t_R \text_out[51]$_DFF_P_  (.CLK(clk),
    .D(n_12317_o_0),
    .QN(_00805_));
 DFFHQNx1_ASAP7_75t_R \text_out[52]$_DFF_P_  (.CLK(clk),
    .D(n_12318_o_0),
    .QN(_00806_));
 DFFHQNx1_ASAP7_75t_R \text_out[53]$_DFF_P_  (.CLK(clk),
    .D(n_12319_o_0),
    .QN(_00807_));
 DFFHQNx1_ASAP7_75t_R \text_out[54]$_DFF_P_  (.CLK(clk),
    .D(n_12320_o_0),
    .QN(_00808_));
 DFFHQNx1_ASAP7_75t_R \text_out[55]$_DFF_P_  (.CLK(clk),
    .D(n_12321_o_0),
    .QN(_00809_));
 DFFHQNx1_ASAP7_75t_R \text_out[56]$_DFF_P_  (.CLK(clk),
    .D(n_12322_o_0),
    .QN(_00834_));
 DFFHQNx1_ASAP7_75t_R \text_out[57]$_DFF_P_  (.CLK(clk),
    .D(n_12323_o_0),
    .QN(_00835_));
 DFFHQNx1_ASAP7_75t_R \text_out[58]$_DFF_P_  (.CLK(clk),
    .D(n_12324_o_0),
    .QN(_00836_));
 DFFHQNx1_ASAP7_75t_R \text_out[59]$_DFF_P_  (.CLK(clk),
    .D(n_12325_o_0),
    .QN(_00837_));
 DFFHQNx1_ASAP7_75t_R \text_out[5]$_DFF_P_  (.CLK(clk),
    .D(n_12351_o_0),
    .QN(_00735_));
 DFFHQNx1_ASAP7_75t_R \text_out[60]$_DFF_P_  (.CLK(clk),
    .D(n_12326_o_0),
    .QN(_00838_));
 DFFHQNx1_ASAP7_75t_R \text_out[61]$_DFF_P_  (.CLK(clk),
    .D(n_12327_o_0),
    .QN(_00839_));
 DFFHQNx1_ASAP7_75t_R \text_out[62]$_DFF_P_  (.CLK(clk),
    .D(n_12328_o_0),
    .QN(_00840_));
 DFFHQNx1_ASAP7_75t_R \text_out[63]$_DFF_P_  (.CLK(clk),
    .D(n_12329_o_0),
    .QN(_00841_));
 DFFHQNx1_ASAP7_75t_R \text_out[64]$_DFF_P_  (.CLK(clk),
    .D(n_12330_o_0),
    .QN(_00746_));
 DFFHQNx1_ASAP7_75t_R \text_out[65]$_DFF_P_  (.CLK(clk),
    .D(n_12331_o_0),
    .QN(_00747_));
 DFFHQNx1_ASAP7_75t_R \text_out[66]$_DFF_P_  (.CLK(clk),
    .D(n_12332_o_0),
    .QN(_00748_));
 DFFHQNx1_ASAP7_75t_R \text_out[67]$_DFF_P_  (.CLK(clk),
    .D(n_12333_o_0),
    .QN(_00749_));
 DFFHQNx1_ASAP7_75t_R \text_out[68]$_DFF_P_  (.CLK(clk),
    .D(n_12334_o_0),
    .QN(_00750_));
 DFFHQNx1_ASAP7_75t_R \text_out[69]$_DFF_P_  (.CLK(clk),
    .D(n_12335_o_0),
    .QN(_00751_));
 DFFHQNx1_ASAP7_75t_R \text_out[6]$_DFF_P_  (.CLK(clk),
    .D(n_12352_o_0),
    .QN(_00736_));
 DFFHQNx1_ASAP7_75t_R \text_out[70]$_DFF_P_  (.CLK(clk),
    .D(n_12336_o_0),
    .QN(_00752_));
 DFFHQNx1_ASAP7_75t_R \text_out[71]$_DFF_P_  (.CLK(clk),
    .D(n_12337_o_0),
    .QN(_00753_));
 DFFHQNx1_ASAP7_75t_R \text_out[72]$_DFF_P_  (.CLK(clk),
    .D(n_12338_o_0),
    .QN(_00778_));
 DFFHQNx1_ASAP7_75t_R \text_out[73]$_DFF_P_  (.CLK(clk),
    .D(n_12339_o_0),
    .QN(_00779_));
 DFFHQNx1_ASAP7_75t_R \text_out[74]$_DFF_P_  (.CLK(clk),
    .D(n_12340_o_0),
    .QN(_00780_));
 DFFHQNx1_ASAP7_75t_R \text_out[75]$_DFF_P_  (.CLK(clk),
    .D(n_12341_o_0),
    .QN(_00781_));
 DFFHQNx1_ASAP7_75t_R \text_out[76]$_DFF_P_  (.CLK(clk),
    .D(n_12342_o_0),
    .QN(_00782_));
 DFFHQNx1_ASAP7_75t_R \text_out[77]$_DFF_P_  (.CLK(clk),
    .D(n_12343_o_0),
    .QN(_00783_));
 DFFHQNx1_ASAP7_75t_R \text_out[78]$_DFF_P_  (.CLK(clk),
    .D(n_12344_o_0),
    .QN(_00784_));
 DFFHQNx1_ASAP7_75t_R \text_out[79]$_DFF_P_  (.CLK(clk),
    .D(n_12345_o_0),
    .QN(_00785_));
 DFFHQNx1_ASAP7_75t_R \text_out[7]$_DFF_P_  (.CLK(clk),
    .D(n_12353_o_0),
    .QN(_00737_));
 DFFHQNx1_ASAP7_75t_R \text_out[80]$_DFF_P_  (.CLK(clk),
    .D(n_12354_o_0),
    .QN(_00810_));
 DFFHQNx1_ASAP7_75t_R \text_out[81]$_DFF_P_  (.CLK(clk),
    .D(n_12355_o_0),
    .QN(_00811_));
 DFFHQNx1_ASAP7_75t_R \text_out[82]$_DFF_P_  (.CLK(clk),
    .D(n_12356_o_0),
    .QN(_00812_));
 DFFHQNx1_ASAP7_75t_R \text_out[83]$_DFF_P_  (.CLK(clk),
    .D(n_12357_o_0),
    .QN(_00813_));
 DFFHQNx1_ASAP7_75t_R \text_out[84]$_DFF_P_  (.CLK(clk),
    .D(n_12358_o_0),
    .QN(_00814_));
 DFFHQNx1_ASAP7_75t_R \text_out[85]$_DFF_P_  (.CLK(clk),
    .D(n_12359_o_0),
    .QN(_00815_));
 DFFHQNx1_ASAP7_75t_R \text_out[86]$_DFF_P_  (.CLK(clk),
    .D(n_12360_o_0),
    .QN(_00816_));
 DFFHQNx1_ASAP7_75t_R \text_out[87]$_DFF_P_  (.CLK(clk),
    .D(n_12361_o_0),
    .QN(_00817_));
 DFFHQNx1_ASAP7_75t_R \text_out[88]$_DFF_P_  (.CLK(clk),
    .D(n_12362_o_0),
    .QN(_00842_));
 DFFHQNx1_ASAP7_75t_R \text_out[89]$_DFF_P_  (.CLK(clk),
    .D(n_12363_o_0),
    .QN(_00843_));
 DFFHQNx1_ASAP7_75t_R \text_out[8]$_DFF_P_  (.CLK(clk),
    .D(n_12274_o_0),
    .QN(_00762_));
 DFFHQNx1_ASAP7_75t_R \text_out[90]$_DFF_P_  (.CLK(clk),
    .D(n_12364_o_0),
    .QN(_00844_));
 DFFHQNx1_ASAP7_75t_R \text_out[91]$_DFF_P_  (.CLK(clk),
    .D(n_12365_o_0),
    .QN(_00845_));
 DFFHQNx1_ASAP7_75t_R \text_out[92]$_DFF_P_  (.CLK(clk),
    .D(n_12366_o_0),
    .QN(_00846_));
 DFFHQNx1_ASAP7_75t_R \text_out[93]$_DFF_P_  (.CLK(clk),
    .D(n_12367_o_0),
    .QN(_00847_));
 DFFHQNx1_ASAP7_75t_R \text_out[94]$_DFF_P_  (.CLK(clk),
    .D(n_12368_o_0),
    .QN(_00848_));
 DFFHQNx1_ASAP7_75t_R \text_out[95]$_DFF_P_  (.CLK(clk),
    .D(n_12369_o_0),
    .QN(_00849_));
 DFFHQNx1_ASAP7_75t_R \text_out[96]$_DFF_P_  (.CLK(clk),
    .D(n_12242_o_0),
    .QN(_00754_));
 DFFHQNx1_ASAP7_75t_R \text_out[97]$_DFF_P_  (.CLK(clk),
    .D(n_12243_o_0),
    .QN(_00755_));
 DFFHQNx1_ASAP7_75t_R \text_out[98]$_DFF_P_  (.CLK(clk),
    .D(n_12244_o_0),
    .QN(_00756_));
 DFFHQNx1_ASAP7_75t_R \text_out[99]$_DFF_P_  (.CLK(clk),
    .D(n_12245_o_0),
    .QN(_00757_));
 DFFHQNx1_ASAP7_75t_R \text_out[9]$_DFF_P_  (.CLK(clk),
    .D(n_12275_o_0),
    .QN(_00763_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/out[24]$_SDFF_PP1_  (.CLK(clk),
    .D(n_12893_o_0),
    .QN(_00446_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/out[25]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12898_o_0),
    .QN(_00447_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/out[26]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12901_o_0),
    .QN(_00448_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/out[27]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12906_o_0),
    .QN(_00449_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/out[28]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12909_o_0),
    .QN(_00450_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/out[29]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12911_o_0),
    .QN(_00451_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/out[30]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12913_o_0),
    .QN(_00452_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/out[31]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12914_o_0),
    .QN(_00453_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/rcnt[0]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12883_o_0),
    .QN(\u0/r0/rcnt_next[0] ));
 DFFHQNx1_ASAP7_75t_R \u0/r0/rcnt[1]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12885_o_0),
    .QN(_11695_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/rcnt[2]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12888_o_0),
    .QN(_00644_));
 DFFHQNx1_ASAP7_75t_R \u0/r0/rcnt[3]$_SDFF_PP0_  (.CLK(clk),
    .D(n_12891_o_0),
    .QN(_00859_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[0]$_DFF_P_  (.CLK(clk),
    .D(n_2631_o_0),
    .QN(_00425_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[10]$_DFF_P_  (.CLK(clk),
    .D(n_2150_o_0),
    .QN(_00424_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[11]$_DFF_P_  (.CLK(clk),
    .D(n_2195_o_0),
    .QN(_00434_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[12]$_DFF_P_  (.CLK(clk),
    .D(n_2238_o_0),
    .QN(_00435_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[13]$_DFF_P_  (.CLK(clk),
    .D(n_2281_o_0),
    .QN(_00436_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[14]$_DFF_P_  (.CLK(clk),
    .D(n_2321_o_0),
    .QN(_00437_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[15]$_DFF_P_  (.CLK(clk),
    .D(n_2363_o_0),
    .QN(_00438_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[16]$_DFF_P_  (.CLK(clk),
    .D(n_1524_o_0),
    .QN(_00439_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[17]$_DFF_P_  (.CLK(clk),
    .D(n_1588_o_0),
    .QN(_00440_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[18]$_DFF_P_  (.CLK(clk),
    .D(n_1640_o_0),
    .QN(_00417_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[19]$_DFF_P_  (.CLK(clk),
    .D(n_1693_o_0),
    .QN(_00441_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[1]$_DFF_P_  (.CLK(clk),
    .D(n_2709_o_0),
    .QN(_00426_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[20]$_DFF_P_  (.CLK(clk),
    .D(n_1733_o_0),
    .QN(_00442_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[21]$_DFF_P_  (.CLK(clk),
    .D(n_1775_o_0),
    .QN(_00443_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[22]$_DFF_P_  (.CLK(clk),
    .D(n_1816_o_0),
    .QN(_00444_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[23]$_DFF_P_  (.CLK(clk),
    .D(n_1857_o_0),
    .QN(_00445_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[24]$_DFF_P_  (.CLK(clk),
    .D(n_1011_o_0),
    .QN(_00988_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[25]$_DFF_P_  (.CLK(clk),
    .D(n_1066_o_0),
    .QN(_00989_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[26]$_DFF_P_  (.CLK(clk),
    .D(n_1118_o_0),
    .QN(_00990_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[27]$_DFF_P_  (.CLK(clk),
    .D(n_1164_o_0),
    .QN(_00991_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[28]$_DFF_P_  (.CLK(clk),
    .D(n_1207_o_0),
    .QN(_00992_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[29]$_DFF_P_  (.CLK(clk),
    .D(n_1253_o_0),
    .QN(_00993_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[2]$_DFF_P_  (.CLK(clk),
    .D(n_2772_o_0),
    .QN(_00423_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[30]$_DFF_P_  (.CLK(clk),
    .D(n_1295_o_0),
    .QN(_00994_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[31]$_DFF_P_  (.CLK(clk),
    .D(n_1338_o_0),
    .QN(_00995_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[3]$_DFF_P_  (.CLK(clk),
    .D(n_2821_o_0),
    .QN(_00427_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[4]$_DFF_P_  (.CLK(clk),
    .D(n_2871_o_0),
    .QN(_00428_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[5]$_DFF_P_  (.CLK(clk),
    .D(n_2916_o_0),
    .QN(_00429_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[6]$_DFF_P_  (.CLK(clk),
    .D(n_2963_o_0),
    .QN(_00430_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[7]$_DFF_P_  (.CLK(clk),
    .D(n_3003_o_0),
    .QN(_00431_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[8]$_DFF_P_  (.CLK(clk),
    .D(n_2030_o_0),
    .QN(_00432_));
 DFFHQNx1_ASAP7_75t_R \u0/subword[9]$_DFF_P_  (.CLK(clk),
    .D(n_2096_o_0),
    .QN(_00433_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[0]$_DFF_P_  (.CLK(clk),
    .D(n_1916_o_0),
    .QN(_00956_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[10]$_DFF_P_  (.CLK(clk),
    .D(net99),
    .QN(_00966_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[11]$_DFF_P_  (.CLK(clk),
    .D(net71),
    .QN(_00967_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[12]$_DFF_P_  (.CLK(clk),
    .D(n_1363_o_0),
    .QN(_00968_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[13]$_DFF_P_  (.CLK(clk),
    .D(n_1426_o_0),
    .QN(_00969_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[14]$_DFF_P_  (.CLK(clk),
    .D(n_1484_o_0),
    .QN(_00970_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[15]$_DFF_P_  (.CLK(clk),
    .D(n_1521_o_0),
    .QN(_00971_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[16]$_DFF_P_  (.CLK(clk),
    .D(n_933_o_0),
    .QN(_00972_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[17]$_DFF_P_  (.CLK(clk),
    .D(n_864_o_0),
    .QN(_00973_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[18]$_DFF_P_  (.CLK(clk),
    .D(n_881_o_0),
    .QN(_00974_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[19]$_DFF_P_  (.CLK(clk),
    .D(n_878_o_0),
    .QN(_00975_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[1]$_DFF_P_  (.CLK(clk),
    .D(n_1941_o_0),
    .QN(_00957_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[20]$_DFF_P_  (.CLK(clk),
    .D(net16),
    .QN(_00976_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[21]$_DFF_P_  (.CLK(clk),
    .D(n_904_o_0),
    .QN(_00977_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[22]$_DFF_P_  (.CLK(clk),
    .D(n_931_o_0),
    .QN(_00978_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[23]$_DFF_P_  (.CLK(clk),
    .D(n_972_o_0),
    .QN(_00979_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[24]$_DFF_P_  (.CLK(clk),
    .D(net102),
    .QN(_00980_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[25]$_DFF_P_  (.CLK(clk),
    .D(net100),
    .QN(_00981_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[26]$_DFF_P_  (.CLK(clk),
    .D(net101),
    .QN(_00982_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[27]$_DFF_P_  (.CLK(clk),
    .D(n_2507_o_0),
    .QN(_00983_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[28]$_DFF_P_  (.CLK(clk),
    .D(n_2527_o_0),
    .QN(_00984_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[29]$_DFF_P_  (.CLK(clk),
    .D(n_2532_o_0),
    .QN(_00985_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[2]$_DFF_P_  (.CLK(clk),
    .D(n_1898_o_0),
    .QN(_00958_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[30]$_DFF_P_  (.CLK(clk),
    .D(n_2384_o_0),
    .QN(_00986_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[31]$_DFF_P_  (.CLK(clk),
    .D(n_2372_o_0),
    .QN(_00987_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[3]$_DFF_P_  (.CLK(clk),
    .D(net33),
    .QN(_00959_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[4]$_DFF_P_  (.CLK(clk),
    .D(net18),
    .QN(_00960_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[5]$_DFF_P_  (.CLK(clk),
    .D(net31),
    .QN(_00961_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[6]$_DFF_P_  (.CLK(clk),
    .D(n_1873_o_0),
    .QN(_00962_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[7]$_DFF_P_  (.CLK(clk),
    .D(n_2027_o_0),
    .QN(_00963_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[8]$_DFF_P_  (.CLK(clk),
    .D(n_1387_o_0),
    .QN(_00964_));
 DFFHQNx1_ASAP7_75t_R \u0/tmp_w[9]$_DFF_P_  (.CLK(clk),
    .D(n_1380_o_0),
    .QN(_00965_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][0]$_DFF_P_  (.CLK(clk),
    .D(n_12371_o_0),
    .QN(_00860_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][10]$_DFF_P_  (.CLK(clk),
    .D(n_12373_o_0),
    .QN(_00870_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][11]$_DFF_P_  (.CLK(clk),
    .D(n_12376_o_0),
    .QN(_00871_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][12]$_DFF_P_  (.CLK(clk),
    .D(n_12379_o_0),
    .QN(_00872_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][13]$_DFF_P_  (.CLK(clk),
    .D(n_12382_o_0),
    .QN(_00873_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][14]$_DFF_P_  (.CLK(clk),
    .D(n_12384_o_0),
    .QN(_00874_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][15]$_DFF_P_  (.CLK(clk),
    .D(n_12386_o_0),
    .QN(_00875_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][16]$_DFF_P_  (.CLK(clk),
    .D(n_12389_o_0),
    .QN(_00876_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][17]$_DFF_P_  (.CLK(clk),
    .D(n_12392_o_0),
    .QN(_00877_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][18]$_DFF_P_  (.CLK(clk),
    .D(n_12394_o_0),
    .QN(_00878_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][19]$_DFF_P_  (.CLK(clk),
    .D(n_12397_o_0),
    .QN(_00879_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][1]$_DFF_P_  (.CLK(clk),
    .D(n_12399_o_0),
    .QN(_00861_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][20]$_DFF_P_  (.CLK(clk),
    .D(n_12402_o_0),
    .QN(_00880_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][21]$_DFF_P_  (.CLK(clk),
    .D(n_12405_o_0),
    .QN(_00881_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][22]$_DFF_P_  (.CLK(clk),
    .D(n_12407_o_0),
    .QN(_00882_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][23]$_DFF_P_  (.CLK(clk),
    .D(n_12409_o_0),
    .QN(_00883_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][24]$_DFF_P_  (.CLK(clk),
    .D(n_12411_o_0),
    .QN(_00884_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][25]$_DFF_P_  (.CLK(clk),
    .D(n_12413_o_0),
    .QN(_00885_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][26]$_DFF_P_  (.CLK(clk),
    .D(n_12415_o_0),
    .QN(_00886_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][27]$_DFF_P_  (.CLK(clk),
    .D(n_12417_o_0),
    .QN(_00887_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][28]$_DFF_P_  (.CLK(clk),
    .D(n_12419_o_0),
    .QN(_00888_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][29]$_DFF_P_  (.CLK(clk),
    .D(n_12422_o_0),
    .QN(_00889_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][2]$_DFF_P_  (.CLK(clk),
    .D(n_12424_o_0),
    .QN(_00862_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][30]$_DFF_P_  (.CLK(clk),
    .D(n_12427_o_0),
    .QN(_00890_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][31]$_DFF_P_  (.CLK(clk),
    .D(n_12429_o_0),
    .QN(_00891_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][3]$_DFF_P_  (.CLK(clk),
    .D(n_12432_o_0),
    .QN(_00863_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][4]$_DFF_P_  (.CLK(clk),
    .D(n_12435_o_0),
    .QN(_00864_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][5]$_DFF_P_  (.CLK(clk),
    .D(n_12438_o_0),
    .QN(_00865_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][6]$_DFF_P_  (.CLK(clk),
    .D(n_12440_o_0),
    .QN(_00866_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][7]$_DFF_P_  (.CLK(clk),
    .D(n_12442_o_0),
    .QN(_00867_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][8]$_DFF_P_  (.CLK(clk),
    .D(n_12444_o_0),
    .QN(_00868_));
 DFFHQNx1_ASAP7_75t_R \u0/w[0][9]$_DFF_P_  (.CLK(clk),
    .D(n_12446_o_0),
    .QN(_00869_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][0]$_DFF_P_  (.CLK(clk),
    .D(n_12448_o_0),
    .QN(_00892_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][10]$_DFF_P_  (.CLK(clk),
    .D(n_12452_o_0),
    .QN(_00902_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][11]$_DFF_P_  (.CLK(clk),
    .D(n_12454_o_0),
    .QN(_00903_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][12]$_DFF_P_  (.CLK(clk),
    .D(n_12457_o_0),
    .QN(_00904_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][13]$_DFF_P_  (.CLK(clk),
    .D(n_12460_o_0),
    .QN(_00905_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][14]$_DFF_P_  (.CLK(clk),
    .D(n_12462_o_0),
    .QN(_00906_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][15]$_DFF_P_  (.CLK(clk),
    .D(n_12465_o_0),
    .QN(_00907_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][16]$_DFF_P_  (.CLK(clk),
    .D(n_12467_o_0),
    .QN(_00908_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][17]$_DFF_P_  (.CLK(clk),
    .D(n_12469_o_0),
    .QN(_00909_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][18]$_DFF_P_  (.CLK(clk),
    .D(n_12472_o_0),
    .QN(_00910_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][19]$_DFF_P_  (.CLK(clk),
    .D(n_12474_o_0),
    .QN(_00911_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][1]$_DFF_P_  (.CLK(clk),
    .D(n_12476_o_0),
    .QN(_00893_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][20]$_DFF_P_  (.CLK(clk),
    .D(n_12479_o_0),
    .QN(_00912_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][21]$_DFF_P_  (.CLK(clk),
    .D(n_12481_o_0),
    .QN(_00913_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][22]$_DFF_P_  (.CLK(clk),
    .D(n_12483_o_0),
    .QN(_00914_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][23]$_DFF_P_  (.CLK(clk),
    .D(n_12485_o_0),
    .QN(_00915_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][24]$_DFF_P_  (.CLK(clk),
    .D(n_12487_o_0),
    .QN(_00916_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][25]$_DFF_P_  (.CLK(clk),
    .D(n_12489_o_0),
    .QN(_00917_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][26]$_DFF_P_  (.CLK(clk),
    .D(n_12491_o_0),
    .QN(_00918_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][27]$_DFF_P_  (.CLK(clk),
    .D(n_12494_o_0),
    .QN(_00919_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][28]$_DFF_P_  (.CLK(clk),
    .D(n_12497_o_0),
    .QN(_00920_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][29]$_DFF_P_  (.CLK(clk),
    .D(n_12500_o_0),
    .QN(_00921_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][2]$_DFF_P_  (.CLK(clk),
    .D(n_12504_o_0),
    .QN(_00894_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][30]$_DFF_P_  (.CLK(clk),
    .D(n_12507_o_0),
    .QN(_00922_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][31]$_DFF_P_  (.CLK(clk),
    .D(n_12509_o_0),
    .QN(_00923_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][3]$_DFF_P_  (.CLK(clk),
    .D(n_12512_o_0),
    .QN(_00895_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][4]$_DFF_P_  (.CLK(clk),
    .D(n_12515_o_0),
    .QN(_00896_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][5]$_DFF_P_  (.CLK(clk),
    .D(n_12518_o_0),
    .QN(_00897_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][6]$_DFF_P_  (.CLK(clk),
    .D(n_12520_o_0),
    .QN(_00898_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][7]$_DFF_P_  (.CLK(clk),
    .D(n_12522_o_0),
    .QN(_00899_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][8]$_DFF_P_  (.CLK(clk),
    .D(n_12524_o_0),
    .QN(_00900_));
 DFFHQNx1_ASAP7_75t_R \u0/w[1][9]$_DFF_P_  (.CLK(clk),
    .D(n_12526_o_0),
    .QN(_00901_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][0]$_DFF_P_  (.CLK(clk),
    .D(n_12529_o_0),
    .QN(_00924_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][10]$_DFF_P_  (.CLK(clk),
    .D(n_12532_o_0),
    .QN(_00934_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][11]$_DFF_P_  (.CLK(clk),
    .D(n_12535_o_0),
    .QN(_00935_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][12]$_DFF_P_  (.CLK(clk),
    .D(n_12538_o_0),
    .QN(_00936_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][13]$_DFF_P_  (.CLK(clk),
    .D(n_12540_o_0),
    .QN(_00937_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][14]$_DFF_P_  (.CLK(clk),
    .D(n_12542_o_0),
    .QN(_00938_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][15]$_DFF_P_  (.CLK(clk),
    .D(n_12544_o_0),
    .QN(_00939_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][16]$_DFF_P_  (.CLK(clk),
    .D(n_12547_o_0),
    .QN(_00940_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][17]$_DFF_P_  (.CLK(clk),
    .D(n_12550_o_0),
    .QN(_00941_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][18]$_DFF_P_  (.CLK(clk),
    .D(n_12553_o_0),
    .QN(_00942_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][19]$_DFF_P_  (.CLK(clk),
    .D(n_12555_o_0),
    .QN(_00943_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][1]$_DFF_P_  (.CLK(clk),
    .D(n_12558_o_0),
    .QN(_00925_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][20]$_DFF_P_  (.CLK(clk),
    .D(n_12561_o_0),
    .QN(_00944_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][21]$_DFF_P_  (.CLK(clk),
    .D(n_12563_o_0),
    .QN(_00945_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][22]$_DFF_P_  (.CLK(clk),
    .D(n_12566_o_0),
    .QN(_00946_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][23]$_DFF_P_  (.CLK(clk),
    .D(n_12568_o_0),
    .QN(_00947_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][24]$_DFF_P_  (.CLK(clk),
    .D(n_12570_o_0),
    .QN(_00948_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][25]$_DFF_P_  (.CLK(clk),
    .D(n_12573_o_0),
    .QN(_00949_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][26]$_DFF_P_  (.CLK(clk),
    .D(n_12576_o_0),
    .QN(_00950_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][27]$_DFF_P_  (.CLK(clk),
    .D(n_12579_o_0),
    .QN(_00951_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][28]$_DFF_P_  (.CLK(clk),
    .D(n_12582_o_0),
    .QN(_00952_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][29]$_DFF_P_  (.CLK(clk),
    .D(n_12585_o_0),
    .QN(_00953_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][2]$_DFF_P_  (.CLK(clk),
    .D(n_12588_o_0),
    .QN(_00926_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][30]$_DFF_P_  (.CLK(clk),
    .D(n_12590_o_0),
    .QN(_00954_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][31]$_DFF_P_  (.CLK(clk),
    .D(n_12593_o_0),
    .QN(_00955_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][3]$_DFF_P_  (.CLK(clk),
    .D(n_12596_o_0),
    .QN(_00927_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][4]$_DFF_P_  (.CLK(clk),
    .D(n_12598_o_0),
    .QN(_00928_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][5]$_DFF_P_  (.CLK(clk),
    .D(n_12601_o_0),
    .QN(_00929_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][6]$_DFF_P_  (.CLK(clk),
    .D(n_12604_o_0),
    .QN(_00930_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][7]$_DFF_P_  (.CLK(clk),
    .D(n_12607_o_0),
    .QN(_00931_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][8]$_DFF_P_  (.CLK(clk),
    .D(n_12610_o_0),
    .QN(_00932_));
 DFFHQNx1_ASAP7_75t_R \u0/w[2][9]$_DFF_P_  (.CLK(clk),
    .D(n_12613_o_0),
    .QN(_00933_));
 assign done = n_12975_o_0;
 assign text_out[0] = n_12976_o_0;
 assign text_out[100] = n_12977_o_0;
 assign text_out[101] = n_12978_o_0;
 assign text_out[102] = n_12979_o_0;
 assign text_out[103] = n_12980_o_0;
 assign text_out[104] = n_12981_o_0;
 assign text_out[105] = n_12982_o_0;
 assign text_out[106] = n_12983_o_0;
 assign text_out[107] = n_12984_o_0;
 assign text_out[108] = n_12985_o_0;
 assign text_out[109] = n_12986_o_0;
 assign text_out[10] = n_12987_o_0;
 assign text_out[110] = n_12988_o_0;
 assign text_out[111] = n_12989_o_0;
 assign text_out[112] = n_12990_o_0;
 assign text_out[113] = n_12991_o_0;
 assign text_out[114] = n_12992_o_0;
 assign text_out[115] = n_12993_o_0;
 assign text_out[116] = n_12994_o_0;
 assign text_out[117] = n_12995_o_0;
 assign text_out[118] = n_12996_o_0;
 assign text_out[119] = n_12997_o_0;
 assign text_out[11] = n_12998_o_0;
 assign text_out[120] = n_12999_o_0;
 assign text_out[121] = n_13000_o_0;
 assign text_out[122] = n_13001_o_0;
 assign text_out[123] = n_13002_o_0;
 assign text_out[124] = n_13003_o_0;
 assign text_out[125] = n_13004_o_0;
 assign text_out[126] = n_13005_o_0;
 assign text_out[127] = n_13006_o_0;
 assign text_out[12] = n_13007_o_0;
 assign text_out[13] = n_13008_o_0;
 assign text_out[14] = n_13009_o_0;
 assign text_out[15] = n_13010_o_0;
 assign text_out[16] = n_13011_o_0;
 assign text_out[17] = n_13012_o_0;
 assign text_out[18] = n_13013_o_0;
 assign text_out[19] = n_13014_o_0;
 assign text_out[1] = n_13015_o_0;
 assign text_out[20] = n_13016_o_0;
 assign text_out[21] = n_13017_o_0;
 assign text_out[22] = n_13018_o_0;
 assign text_out[23] = n_13019_o_0;
 assign text_out[24] = n_13020_o_0;
 assign text_out[25] = n_13021_o_0;
 assign text_out[26] = n_13022_o_0;
 assign text_out[27] = n_13023_o_0;
 assign text_out[28] = n_13024_o_0;
 assign text_out[29] = n_13025_o_0;
 assign text_out[2] = n_13026_o_0;
 assign text_out[30] = n_13027_o_0;
 assign text_out[31] = n_13028_o_0;
 assign text_out[32] = n_13029_o_0;
 assign text_out[33] = n_13030_o_0;
 assign text_out[34] = n_13031_o_0;
 assign text_out[35] = n_13032_o_0;
 assign text_out[36] = n_13033_o_0;
 assign text_out[37] = n_13034_o_0;
 assign text_out[38] = n_13035_o_0;
 assign text_out[39] = n_13036_o_0;
 assign text_out[3] = n_13037_o_0;
 assign text_out[40] = n_13038_o_0;
 assign text_out[41] = n_13039_o_0;
 assign text_out[42] = n_13040_o_0;
 assign text_out[43] = n_13041_o_0;
 assign text_out[44] = n_13042_o_0;
 assign text_out[45] = n_13043_o_0;
 assign text_out[46] = n_13044_o_0;
 assign text_out[47] = n_13045_o_0;
 assign text_out[48] = n_13046_o_0;
 assign text_out[49] = n_13047_o_0;
 assign text_out[4] = n_13048_o_0;
 assign text_out[50] = n_13049_o_0;
 assign text_out[51] = n_13050_o_0;
 assign text_out[52] = n_13051_o_0;
 assign text_out[53] = n_13052_o_0;
 assign text_out[54] = n_13053_o_0;
 assign text_out[55] = n_13054_o_0;
 assign text_out[56] = n_13055_o_0;
 assign text_out[57] = n_13056_o_0;
 assign text_out[58] = n_13057_o_0;
 assign text_out[59] = n_13058_o_0;
 assign text_out[5] = n_13059_o_0;
 assign text_out[60] = n_13060_o_0;
 assign text_out[61] = n_13061_o_0;
 assign text_out[62] = n_13062_o_0;
 assign text_out[63] = n_13063_o_0;
 assign text_out[64] = n_13064_o_0;
 assign text_out[65] = n_13065_o_0;
 assign text_out[66] = n_13066_o_0;
 assign text_out[67] = n_13067_o_0;
 assign text_out[68] = n_13068_o_0;
 assign text_out[69] = n_13069_o_0;
 assign text_out[6] = n_13070_o_0;
 assign text_out[70] = n_13071_o_0;
 assign text_out[71] = n_13072_o_0;
 assign text_out[72] = n_13073_o_0;
 assign text_out[73] = n_13074_o_0;
 assign text_out[74] = n_13075_o_0;
 assign text_out[75] = n_13076_o_0;
 assign text_out[76] = n_13077_o_0;
 assign text_out[77] = n_13078_o_0;
 assign text_out[78] = n_13079_o_0;
 assign text_out[79] = n_13080_o_0;
 assign text_out[7] = n_13081_o_0;
 assign text_out[80] = n_13082_o_0;
 assign text_out[81] = n_13083_o_0;
 assign text_out[82] = n_13084_o_0;
 assign text_out[83] = n_13085_o_0;
 assign text_out[84] = n_13086_o_0;
 assign text_out[85] = n_13087_o_0;
 assign text_out[86] = n_13088_o_0;
 assign text_out[87] = n_13089_o_0;
 assign text_out[88] = n_13090_o_0;
 assign text_out[89] = n_13091_o_0;
 assign text_out[8] = n_13092_o_0;
 assign text_out[90] = n_13093_o_0;
 assign text_out[91] = n_13094_o_0;
 assign text_out[92] = n_13095_o_0;
 assign text_out[93] = n_13096_o_0;
 assign text_out[94] = n_13097_o_0;
 assign text_out[95] = n_13098_o_0;
 assign text_out[96] = n_13099_o_0;
 assign text_out[97] = n_13100_o_0;
 assign text_out[98] = n_13101_o_0;
 assign text_out[99] = n_13102_o_0;
 assign text_out[9] = n_13103_o_0;
endmodule
